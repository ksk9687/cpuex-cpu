library IEEE;
use IEEE.std_logic_1164.all;

library work;

package fp_inv_table is

subtype vec24 is std_logic_vector(23 downto 0);
type table_t is array (0 to 2047) of vec24;
constant table : table_t := (
"111111111110000000000010",
"111111111010000000011010",
"111111110110000001001010",
"111111110010000010010010",
"111111101110000011110010",
"111111101010000101101001",
"111111100110000111111000",
"111111100010001010011111",
"111111011110001101011110",
"111111011010010000110100",
"111111010110010100100010",
"111111010010011000100111",
"111111001110011101000011",
"111111001010100001110111",
"111111000110100111000011",
"111111000010101100100110",
"111110111110110010100000",
"111110111010111000110001",
"111110110110111111011010",
"111110110011000110011001",
"111110101111001101110000",
"111110101011010101011110",
"111110100111011101100011",
"111110100011100101111111",
"111110011111101110110001",
"111110011011110111111011",
"111110011000000001011011",
"111110010100001011010011",
"111110010000010101100001",
"111110001100100000000101",
"111110001000101011000001",
"111110000100110110010011",
"111110000001000001111100",
"111101111101001101111011",
"111101111001011010010000",
"111101110101100110111100",
"111101110001110011111111",
"111101101110000001011000",
"111101101010001111000111",
"111101100110011101001100",
"111101100010101011101000",
"111101011110111010011010",
"111101011011001001100010",
"111101010111011001000000",
"111101010011101000110100",
"111101001111111000111110",
"111101001100001001011111",
"111101001000011010010101",
"111101000100101011100001",
"111101000000111101000011",
"111100111101001110111010",
"111100111001100001001000",
"111100110101110011101011",
"111100110010000110100100",
"111100101110011001110011",
"111100101010101101010111",
"111100100111000001010000",
"111100100011010101100000",
"111100011111101010000100",
"111100011011111110111111",
"111100011000010100001110",
"111100010100101001110011",
"111100010000111111101101",
"111100001101010101111101",
"111100001001101100100010",
"111100000110000011011100",
"111100000010011010101011",
"111011111110110010001111",
"111011111011001010001000",
"111011110111100010010111",
"111011110011111010111010",
"111011110000010011110010",
"111011101100101101000000",
"111011101001000110100010",
"111011100101100000011001",
"111011100001111010100101",
"111011011110010101000101",
"111011011010101111111010",
"111011010111001011000100",
"111011010011100110100011",
"111011010000000010010110",
"111011001100011110011110",
"111011001000111010111010",
"111011000101010111101011",
"111011000001110100110000",
"111010111110010010001010",
"111010111010101111111000",
"111010110111001101111011",
"111010110011101100010001",
"111010110000001010111100",
"111010101100101001111011",
"111010101001001001001111",
"111010100101101000110110",
"111010100010001000110010",
"111010011110101001000010",
"111010011011001001100110",
"111010010111101010011101",
"111010010100001011101001",
"111010010000101101001001",
"111010001101001110111100",
"111010001001110001000100",
"111010000110010011011111",
"111010000010110110001110",
"111001111111011001010000",
"111001111011111100100111",
"111001111000100000010001",
"111001110101000100001111",
"111001110001101000100000",
"111001101110001101000101",
"111001101010110001111101",
"111001100111010111001001",
"111001100011111100101001",
"111001100000100010011011",
"111001011101001000100001",
"111001011001101110111011",
"111001010110010101101000",
"111001010010111100101000",
"111001001111100011111011",
"111001001100001011100010",
"111001001000110011011011",
"111001000101011011101000",
"111001000010000100001000",
"111000111110101100111011",
"111000111011010110000001",
"111000110111111111011010",
"111000110100101001000110",
"111000110001010011000100",
"111000101101111101010110",
"111000101010100111111011",
"111000100111010010110010",
"111000100011111101111100",
"111000100000101001011001",
"111000011101010101001001",
"111000011010000001001011",
"111000010110101101100000",
"111000010011011010000111",
"111000010000000111000010",
"111000001100110100001110",
"111000001001100001101101",
"111000000110001111011111",
"111000000010111101100011",
"110111111111101011111001",
"110111111100011010100010",
"110111111001001001011101",
"110111110101111000101011",
"110111110010101000001011",
"110111101111010111111101",
"110111101100001000000001",
"110111101000111000010111",
"110111100101101001000000",
"110111100010011001111010",
"110111011111001011000111",
"110111011011111100100110",
"110111011000101110010111",
"110111010101100000011001",
"110111010010010010101110",
"110111001111000101010101",
"110111001011111000001101",
"110111001000101011010111",
"110111000101011110110011",
"110111000010010010100001",
"110110111111000110100001",
"110110111011111010110010",
"110110111000101111010101",
"110110110101100100001010",
"110110110010011001010000",
"110110101111001110101000",
"110110101100000100010001",
"110110101000111010001100",
"110110100101110000011001",
"110110100010100110110111",
"110110011111011101100110",
"110110011100010100100111",
"110110011001001011111001",
"110110010110000011011100",
"110110010010111011010001",
"110110001111110011010111",
"110110001100101011101110",
"110110001001100100010111",
"110110000110011101010001",
"110110000011010110011011",
"110110000000001111110111",
"110101111101001001100100",
"110101111010000011100010",
"110101110110111101110010",
"110101110011111000010010",
"110101110000110011000011",
"110101101101101110000101",
"110101101010101001011000",
"110101100111100100111011",
"110101100100100000110000",
"110101100001011100110101",
"110101011110011001001100",
"110101011011010101110011",
"110101011000010010101010",
"110101010101001111110011",
"110101010010001101001100",
"110101001111001010110110",
"110101001100001000110000",
"110101001001000110111011",
"110101000110000101010110",
"110101000011000100000010",
"110101000000000010111111",
"110100111101000010001100",
"110100111010000001101001",
"110100110111000001010111",
"110100110100000001010101",
"110100110001000001100011",
"110100101110000010000010",
"110100101011000010110001",
"110100101000000011110000",
"110100100101000101000000",
"110100100010000110100000",
"110100011111001000001111",
"110100011100001010001111",
"110100011001001100100000",
"110100010110001111000000",
"110100010011010001110000",
"110100010000010100110001",
"110100001101011000000001",
"110100001010011011100001",
"110100000111011111010001",
"110100000100100011010010",
"110100000001100111100010",
"110011111110101100000001",
"110011111011110000110001",
"110011111000110101110001",
"110011110101111011000000",
"110011110011000000011111",
"110011110000000110001110",
"110011101101001100001100",
"110011101010010010011010",
"110011100111011000111000",
"110011100100011111100110",
"110011100001100110100011",
"110011011110101101101111",
"110011011011110101001011",
"110011011000111100110111",
"110011010110000100110010",
"110011010011001100111100",
"110011010000010101010110",
"110011001101011101111111",
"110011001010100110111000",
"110011000111110000000000",
"110011000100111001010111",
"110011000010000010111110",
"110010111111001100110100",
"110010111100010110111001",
"110010111001100001001101",
"110010110110101011110001",
"110010110011110110100011",
"110010110001000001100101",
"110010101110001100110110",
"110010101011011000010110",
"110010101000100100000101",
"110010100101110000000011",
"110010100010111100010000",
"110010100000001000101100",
"110010011101010101010111",
"110010011010100010010000",
"110010010111101111011001",
"110010010100111100110001",
"110010010010001010010111",
"110010001111011000001100",
"110010001100100110010000",
"110010001001110100100011",
"110010000111000011000101",
"110010000100010001110101",
"110010000001100000110100",
"110001111110110000000010",
"110001111011111111011110",
"110001111001001111001001",
"110001110110011111000010",
"110001110011101111001010",
"110001110000111111100001",
"110001101110010000000110",
"110001101011100000111001",
"110001101000110001111011",
"110001100110000011001100",
"110001100011010100101010",
"110001100000100110011000",
"110001011101111000010011",
"110001011011001010011101",
"110001011000011100110101",
"110001010101101111011100",
"110001010011000010010001",
"110001010000010101010100",
"110001001101101000100101",
"110001001010111100000100",
"110001001000001111110010",
"110001000101100011101110",
"110001000010110111111000",
"110001000000001100010000",
"110000111101100000110110",
"110000111010110101101010",
"110000111000001010101100",
"110000110101011111111100",
"110000110010110101011010",
"110000110000001011000110",
"110000101101100001000000",
"110000101010110111001000",
"110000101000001101011101",
"110000100101100100000001",
"110000100010111010110010",
"110000100000010001110010",
"110000011101101000111111",
"110000011011000000011001",
"110000011000011000000010",
"110000010101101111111000",
"110000010011000111111100",
"110000010000100000001110",
"110000001101111000101101",
"110000001011010001011010",
"110000001000101010010100",
"110000000110000011011100",
"110000000011011100110010",
"110000000000110110010101",
"101111111110010000000110",
"101111111011101010000100",
"101111111001000100001111",
"101111110110011110101000",
"101111110011111001001111",
"101111110001010100000010",
"101111101110101111000100",
"101111101100001010010010",
"101111101001100101101110",
"101111100111000001010111",
"101111100100011101001110",
"101111100001111001010001",
"101111011111010101100010",
"101111011100110010000000",
"101111011010001110101100",
"101111010111101011100100",
"101111010101001000101010",
"101111010010100101111101",
"101111010000000011011101",
"101111001101100001001010",
"101111001010111111000100",
"101111001000011101001011",
"101111000101111011011111",
"101111000011011010000000",
"101111000000111000101110",
"101110111110010111101001",
"101110111011110110110001",
"101110111001010110000110",
"101110110110110101100111",
"101110110100010101010110",
"101110110001110101010010",
"101110101111010101011010",
"101110101100110101101111",
"101110101010010110010001",
"101110100111110110111111",
"101110100101010111111011",
"101110100010111001000011",
"101110100000011010010111",
"101110011101111011111001",
"101110011011011101100111",
"101110011000111111100010",
"101110010110100001101001",
"101110010100000011111101",
"101110010001100110011101",
"101110001111001001001010",
"101110001100101100000100",
"101110001010001111001010",
"101110000111110010011100",
"101110000101010101111011",
"101110000010111001100111",
"101110000000011101011111",
"101101111110000001100011",
"101101111011100101110100",
"101101111001001010010001",
"101101110110101110111010",
"101101110100010011110000",
"101101110001111000110010",
"101101101111011110000000",
"101101101101000011011010",
"101101101010101001000001",
"101101101000001110110100",
"101101100101110100110011",
"101101100011011010111111",
"101101100001000001010110",
"101101011110100111111010",
"101101011100001110101010",
"101101011001110101100101",
"101101010111011100101101",
"101101010101000100000001",
"101101010010101011100001",
"101101010000010011001101",
"101101001101111011000101",
"101101001011100011001010",
"101101001001001011011010",
"101101000110110011110101",
"101101000100011100011101",
"101101000010000101010001",
"101100111111101110010001",
"101100111101010111011100",
"101100111011000000110100",
"101100111000101010010111",
"101100110110010100000110",
"101100110011111110000000",
"101100110001101000000111",
"101100101111010010011001",
"101100101100111100110111",
"101100101010100111100001",
"101100101000010010010110",
"101100100101111101011000",
"101100100011101000100100",
"101100100001010011111101",
"101100011110111111100001",
"101100011100101011010000",
"101100011010010111001011",
"101100011000000011010010",
"101100010101101111100100",
"101100010011011100000010",
"101100010001001000101011",
"101100001110110101100000",
"101100001100100010100000",
"101100001010001111101100",
"101100000111111101000011",
"101100000101101010100101",
"101100000011011000010011",
"101100000001000110001101",
"101011111110110100010001",
"101011111100100010100001",
"101011111010010000111100",
"101011110111111111100011",
"101011110101101110010101",
"101011110011011101010010",
"101011110001001100011010",
"101011101110111011101110",
"101011101100101011001100",
"101011101010011010110110",
"101011101000001010101100",
"101011100101111010101100",
"101011100011101010110111",
"101011100001011011001110",
"101011011111001011101111",
"101011011100111100011100",
"101011011010101101010100",
"101011011000011110010111",
"101011010110001111100100",
"101011010100000000111101",
"101011010001110010100001",
"101011001111100100010000",
"101011001101010110001010",
"101011001011001000001110",
"101011001000111010011110",
"101011000110101100111001",
"101011000100011111011110",
"101011000010010010001110",
"101011000000000101001010",
"101010111101111000010000",
"101010111011101011100000",
"101010111001011110111100",
"101010110111010010100010",
"101010110101000110010011",
"101010110010111010001111",
"101010110000101110010110",
"101010101110100010100111",
"101010101100010111000011",
"101010101010001011101010",
"101010101000000000011011",
"101010100101110101010111",
"101010100011101010011110",
"101010100001011111101111",
"101010011111010101001011",
"101010011101001010110010",
"101010011011000000100011",
"101010011000110110011110",
"101010010110101100100100",
"101010010100100010110101",
"101010010010011001010000",
"101010010000001111110110",
"101010001110000110100110",
"101010001011111101100000",
"101010001001110100100101",
"101010000111101011110100",
"101010000101100011001110",
"101010000011011010110010",
"101010000001010010100000",
"101001111111001010011001",
"101001111101000010011100",
"101001111010111010101010",
"101001111000110011000010",
"101001110110101011100100",
"101001110100100100010000",
"101001110010011101000110",
"101001110000010110000111",
"101001101110001111010010",
"101001101100001000100111",
"101001101010000010000111",
"101001100111111011110000",
"101001100101110101100100",
"101001100011101111100010",
"101001100001101001101001",
"101001011111100011111100",
"101001011101011110011000",
"101001011011011000111110",
"101001011001010011101110",
"101001010111001110101000",
"101001010101001001101101",
"101001010011000100111011",
"101001010001000000010011",
"101001001110111011110110",
"101001001100110111100010",
"101001001010110011011000",
"101001001000101111011000",
"101001000110101011100010",
"101001000100100111110110",
"101001000010100100010100",
"101001000000100000111100",
"101000111110011101101101",
"101000111100011010101001",
"101000111010010111101110",
"101000111000010100111101",
"101000110110010010010110",
"101000110100001111111000",
"101000110010001101100101",
"101000110000001011011011",
"101000101110001001011011",
"101000101100000111100100",
"101000101010000101110111",
"101000101000000100010100",
"101000100110000010111011",
"101000100100000001101011",
"101000100010000000100101",
"101000011111111111101001",
"101000011101111110110110",
"101000011011111110001100",
"101000011001111101101101",
"101000010111111101010111",
"101000010101111101001010",
"101000010011111101000111",
"101000010001111101001110",
"101000001111111101011110",
"101000001101111101110111",
"101000001011111110011010",
"101000001001111111000110",
"101000000111111111111100",
"101000000110000000111100",
"101000000100000010000100",
"101000000010000011010110",
"101000000000000100110010",
"100111111110000110010111",
"100111111100001000000101",
"100111111010001001111101",
"100111111000001011111110",
"100111110110001110001000",
"100111110100010000011100",
"100111110010010010111000",
"100111110000010101011110",
"100111101110011000001110",
"100111101100011011000111",
"100111101010011110001000",
"100111101000100001010011",
"100111100110100100101000",
"100111100100101000000101",
"100111100010101011101100",
"100111100000101111011100",
"100111011110110011010101",
"100111011100110111010111",
"100111011010111011100010",
"100111011000111111110110",
"100111010111000100010100",
"100111010101001000111010",
"100111010011001101101010",
"100111010001010010100010",
"100111001111010111100100",
"100111001101011100101111",
"100111001011100010000010",
"100111001001100111011111",
"100111000111101101000101",
"100111000101110010110011",
"100111000011111000101011",
"100111000001111110101011",
"100111000000000100110101",
"100110111110001011000111",
"100110111100010001100010",
"100110111010011000000110",
"100110111000011110110011",
"100110110110100101101001",
"100110110100101100101000",
"100110110010110011110000",
"100110110000111011000000",
"100110101111000010011001",
"100110101101001001111011",
"100110101011010001100110",
"100110101001011001011001",
"100110100111100001010101",
"100110100101101001011010",
"100110100011110001101000",
"100110100001111001111111",
"100110100000000010011110",
"100110011110001011000101",
"100110011100010011110110",
"100110011010011100101111",
"100110011000100101110001",
"100110010110101110111011",
"100110010100111000001110",
"100110010011000001101010",
"100110010001001011001110",
"100110001111010100111011",
"100110001101011110110000",
"100110001011101000101110",
"100110001001110010110101",
"100110000111111101000100",
"100110000110000111011011",
"100110000100010001111011",
"100110000010011100100100",
"100110000000100111010101",
"100101111110110010001110",
"100101111100111101010000",
"100101111011001000011011",
"100101111001010011101101",
"100101110111011111001001",
"100101110101101010101100",
"100101110011110110011000",
"100101110010000010001100",
"100101110000001110001001",
"100101101110011010001110",
"100101101100100110011100",
"100101101010110010110001",
"100101101000111111010000",
"100101100111001011110110",
"100101100101011000100101",
"100101100011100101011011",
"100101100001110010011011",
"100101011111111111100010",
"100101011110001100110010",
"100101011100011010001010",
"100101011010100111101010",
"100101011000110101010010",
"100101010111000011000011",
"100101010101010000111011",
"100101010011011110111100",
"100101010001101101000101",
"100101001111111011010110",
"100101001110001001110000",
"100101001100011000010001",
"100101001010100110111011",
"100101001000110101101100",
"100101000111000100100110",
"100101000101010011101000",
"100101000011100010110001",
"100101000001110010000011",
"100101000000000001011101",
"100100111110010000111111",
"100100111100100000101001",
"100100111010110000011011",
"100100111001000000010101",
"100100110111010000010111",
"100100110101100000100001",
"100100110011110000110010",
"100100110010000001001100",
"100100110000010001101110",
"100100101110100010010111",
"100100101100110011001001",
"100100101011000100000010",
"100100101001010101000011",
"100100100111100110001101",
"100100100101110111011110",
"100100100100001000110110",
"100100100010011010010111",
"100100100000101011111111",
"100100011110111101110000",
"100100011101001111101000",
"100100011011100001101000",
"100100011001110011101111",
"100100011000000101111111",
"100100010110011000010110",
"100100010100101010110101",
"100100010010111101011100",
"100100010001010000001010",
"100100001111100011000000",
"100100001101110101111110",
"100100001100001001000011",
"100100001010011100010000",
"100100001000101111100101",
"100100000111000011000010",
"100100000101010110100110",
"100100000011101010010001",
"100100000001111110000101",
"100100000000010010000000",
"100011111110100110000010",
"100011111100111010001100",
"100011111011001110011110",
"100011111001100010110111",
"100011110111110111011000",
"100011110110001100000000",
"100011110100100000110000",
"100011110010110101101000",
"100011110001001010100110",
"100011101111011111101101",
"100011101101110100111011",
"100011101100001010010000",
"100011101010011111101101",
"100011101000110101010001",
"100011100111001010111101",
"100011100101100000110000",
"100011100011110110101011",
"100011100010001100101101",
"100011100000100010110110",
"100011011110111001000111",
"100011011101001111011111",
"100011011011100101111110",
"100011011001111100100101",
"100011011000010011010011",
"100011010110101010001001",
"100011010101000001000110",
"100011010011011000001010",
"100011010001101111010101",
"100011010000000110101000",
"100011001110011110000010",
"100011001100110101100100",
"100011001011001101001100",
"100011001001100100111100",
"100011000111111100110011",
"100011000110010100110001",
"100011000100101100110111",
"100011000011000101000100",
"100011000001011101011000",
"100010111111110101110011",
"100010111110001110010101",
"100010111100100110111110",
"100010111010111111101111",
"100010111001011000100111",
"100010110111110001100110",
"100010110110001010101100",
"100010110100100011111001",
"100010110010111101001101",
"100010110001010110101000",
"100010101111110000001011",
"100010101110001001110100",
"100010101100100011100101",
"100010101010111101011100",
"100010101001010111011011",
"100010100111110001100001",
"100010100110001011101101",
"100010100100100110000001",
"100010100011000000011100",
"100010100001011010111110",
"100010011111110101100110",
"100010011110010000010110",
"100010011100101011001101",
"100010011011000110001010",
"100010011001100001001111",
"100010010111111100011010",
"100010010110010111101100",
"100010010100110011000110",
"100010010011001110100110",
"100010010001101010001101",
"100010010000000101111011",
"100010001110100001110000",
"100010001100111101101100",
"100010001011011001101110",
"100010001001110101111000",
"100010001000010010001000",
"100010000110101110011111",
"100010000101001010111101",
"100010000011100111100010",
"100010000010000100001101",
"100010000000100000111111",
"100001111110111101111000",
"100001111101011010111000",
"100001111011110111111111",
"100001111010010101001100",
"100001111000110010100000",
"100001110111001111111011",
"100001110101101101011100",
"100001110100001011000101",
"100001110010101000110100",
"100001110001000110101001",
"100001101111100100100110",
"100001101110000010101000",
"100001101100100000110010",
"100001101010111111000010",
"100001101001011101011001",
"100001100111111011110111",
"100001100110011010011011",
"100001100100111001000110",
"100001100011010111110111",
"100001100001110110101111",
"100001100000010101101110",
"100001011110110100110011",
"100001011101010011111111",
"100001011011110011010001",
"100001011010010010101010",
"100001011000110010001001",
"100001010111010001101111",
"100001010101110001011100",
"100001010100010001001111",
"100001010010110001001000",
"100001010001010001001000",
"100001001111110001001110",
"100001001110010001011011",
"100001001100110001101111",
"100001001011010010001001",
"100001001001110010101001",
"100001001000010011010000",
"100001000110110011111101",
"100001000101010100110000",
"100001000011110101101010",
"100001000010010110101011",
"100001000000110111110001",
"100000111111011000111111",
"100000111101111010010010",
"100000111100011011101100",
"100000111010111101001100",
"100000111001011110110011",
"100000111000000000100000",
"100000110110100010010011",
"100000110101000100001101",
"100000110011100110001101",
"100000110010001000010011",
"100000110000101010100000",
"100000101111001100110011",
"100000101101101111001100",
"100000101100010001101011",
"100000101010110100010001",
"100000101001010110111101",
"100000100111111001101111",
"100000100110011100100111",
"100000100100111111100110",
"100000100011100010101011",
"100000100010000101110110",
"100000100000101001000111",
"100000011111001100011110",
"100000011101101111111100",
"100000011100010011100000",
"100000011010110111001010",
"100000011001011010111010",
"100000010111111110110000",
"100000010110100010101100",
"100000010101000110101111",
"100000010011101010111000",
"100000010010001111000110",
"100000010000110011011011",
"100000001111010111110110",
"100000001101111100010111",
"100000001100100000111111",
"100000001011000101101100",
"100000001001101010011111",
"100000001000001111011001",
"100000000110110100011000",
"100000000101011001011101",
"100000000011111110101001",
"100000000010100011111010",
"100000000001001001010010",
"011111111111101110101111",
"011111111110010100010011",
"011111111100111001111100",
"011111111011011111101100",
"011111111010000101100001",
"011111111000101011011101",
"011111110111010001011110",
"011111110101110111100110",
"011111110100011101110011",
"011111110011000100000110",
"011111110001101010011111",
"011111110000010000111110",
"011111101110110111100011",
"011111101101011110001110",
"011111101100000100111111",
"011111101010101011110101",
"011111101001010010110010",
"011111100111111001110100",
"011111100110100000111101",
"011111100101001000001011",
"011111100011101111011111",
"011111100010010110111000",
"011111100000111110011000",
"011111011111100101111101",
"011111011110001101101001",
"011111011100110101011010",
"011111011011011101010001",
"011111011010000101001101",
"011111011000101101010000",
"011111010111010101011000",
"011111010101111101100110",
"011111010100100101111001",
"011111010011001110010011",
"011111010001110110110010",
"011111010000011111010111",
"011111001111001000000001",
"011111001101110000110010",
"011111001100011001101000",
"011111001011000010100100",
"011111001001101011100101",
"011111001000010100101100",
"011111000110111101111001",
"011111000101100111001100",
"011111000100010000100100",
"011111000010111010000010",
"011111000001100011100101",
"011111000000001101001110",
"011110111110110110111101",
"011110111101100000110001",
"011110111100001010101011",
"011110111010110100101011",
"011110111001011110110000",
"011110111000001000111011",
"011110110110110011001011",
"011110110101011101100001",
"011110110100000111111101",
"011110110010110010011110",
"011110110001011101000100",
"011110110000000111110000",
"011110101110110010100010",
"011110101101011101011001",
"011110101100001000010110",
"011110101010110011011000",
"011110101001011110100000",
"011110101000001001101110",
"011110100110110101000000",
"011110100101100000011001",
"011110100100001011110110",
"011110100010110111011010",
"011110100001100011000010",
"011110100000001110110001",
"011110011110111010100100",
"011110011101100110011101",
"011110011100010010011100",
"011110011010111110100000",
"011110011001101010101001",
"011110011000010110111000",
"011110010111000011001100",
"011110010101101111100110",
"011110010100011100000101",
"011110010011001000101001",
"011110010001110101010011",
"011110010000100010000010",
"011110001111001110110110",
"011110001101111011110000",
"011110001100101000101111",
"011110001011010101110100",
"011110001010000010111110",
"011110001000110000001101",
"011110000111011101100010",
"011110000110001010111011",
"011110000100111000011011",
"011110000011100101111111",
"011110000010010011101001",
"011110000001000001011000",
"011101111111101111001100",
"011101111110011101000110",
"011101111101001011000101",
"011101111011111001001001",
"011101111010100111010010",
"011101111001010101100001",
"011101111000000011110100",
"011101110110110010001101",
"011101110101100000101100",
"011101110100001111001111",
"011101110010111101111000",
"011101110001101100100110",
"011101110000011011011001",
"011101101111001010010001",
"011101101101111001001111",
"011101101100101000010001",
"011101101011010111011001",
"011101101010000110100110",
"011101101000110101111000",
"011101100111100101010000",
"011101100110010100101100",
"011101100101000100001110",
"011101100011110011110100",
"011101100010100011100000",
"011101100001010011010001",
"011101100000000011000111",
"011101011110110011000010",
"011101011101100011000010",
"011101011100010011001000",
"011101011011000011010010",
"011101011001110011100001",
"011101011000100011110110",
"011101010111010100010000",
"011101010110000100101110",
"011101010100110101010010",
"011101010011100101111011",
"011101010010010110101000",
"011101010001000111011011",
"011101001111111000010011",
"011101001110101001010000",
"011101001101011010010001",
"011101001100001011011000",
"011101001010111100100100",
"011101001001101101110101",
"011101001000011111001011",
"011101000111010000100101",
"011101000110000010000101",
"011101000100110011101010",
"011101000011100101010011",
"011101000010010111000010",
"011101000001001000110101",
"011100111111111010101110",
"011100111110101100101011",
"011100111101011110101101",
"011100111100010000110101",
"011100111011000011000001",
"011100111001110101010010",
"011100111000100111101000",
"011100110111011010000010",
"011100110110001100100010",
"011100110100111111000111",
"011100110011110001110000",
"011100110010100100011110",
"011100110001010111010001",
"011100110000001010001001",
"011100101110111101000110",
"011100101101110000001000",
"011100101100100011001110",
"011100101011010110011010",
"011100101010001001101010",
"011100101000111100111111",
"011100100111110000011001",
"011100100110100011110111",
"011100100101010111011011",
"011100100100001011000011",
"011100100010111110110000",
"011100100001110010100001",
"011100100000100110011000",
"011100011111011010010011",
"011100011110001110010011",
"011100011101000010011000",
"011100011011110110100001",
"011100011010101010101111",
"011100011001011111000010",
"011100011000010011011010",
"011100010111000111110111",
"011100010101111100011000",
"011100010100110000111101",
"011100010011100101101000",
"011100010010011010010111",
"011100010001001111001011",
"011100010000000100000100",
"011100001110111001000001",
"011100001101101110000011",
"011100001100100011001001",
"011100001011011000010101",
"011100001010001101100101",
"011100001001000010111001",
"011100000111111000010010",
"011100000110101101110000",
"011100000101100011010011",
"011100000100011000111010",
"011100000011001110100101",
"011100000010000100010110",
"011100000000111010001011",
"011011111111110000000100",
"011011111110100110000010",
"011011111101011100000101",
"011011111100010010001100",
"011011111011001000011000",
"011011111001111110101000",
"011011111000110100111101",
"011011110111101011010111",
"011011110110100001110101",
"011011110101011000011000",
"011011110100001110111111",
"011011110011000101101010",
"011011110001111100011011",
"011011110000110011001111",
"011011101111101010001001",
"011011101110100001000110",
"011011101101011000001001",
"011011101100001111001111",
"011011101011000110011011",
"011011101001111101101011",
"011011101000110100111111",
"011011100111101100010111",
"011011100110100011110101",
"011011100101011011010110",
"011011100100010010111100",
"011011100011001010100111",
"011011100010000010010110",
"011011100000111010001001",
"011011011111110010000001",
"011011011110101001111110",
"011011011101100001111110",
"011011011100011010000100",
"011011011011010010001101",
"011011011010001010011011",
"011011011001000010101101",
"011011010111111011000100",
"011011010110110011011111",
"011011010101101011111111",
"011011010100100100100011",
"011011010011011101001011",
"011011010010010101111000",
"011011010001001110101001",
"011011010000000111011110",
"011011001111000000011000",
"011011001101111001010110",
"011011001100110010011001",
"011011001011101011011111",
"011011001010100100101010",
"011011001001011101111010",
"011011001000010111001110",
"011011000111010000100110",
"011011000110001010000010",
"011011000101000011100011",
"011011000011111101001000",
"011011000010110110110001",
"011011000001110000011110",
"011011000000101010010000",
"011010111111100100000110",
"011010111110011110000001",
"011010111101010111111111",
"011010111100010010000010",
"011010111011001100001001",
"011010111010000110010101",
"011010111001000000100100",
"011010110111111010111000",
"011010110110110101010000",
"011010110101101111101100",
"011010110100101010001101",
"011010110011100100110010",
"011010110010011111011011",
"011010110001011010001000",
"011010110000010100111001",
"011010101111001111101111",
"011010101110001010101001",
"011010101101000101100111",
"011010101100000000101001",
"011010101010111011101111",
"011010101001110110111001",
"011010101000110010001000",
"011010100111101101011011",
"011010100110101000110010",
"011010100101100100001101",
"011010100100011111101100",
"011010100011011011001111",
"011010100010010110110111",
"011010100001010010100010",
"011010100000001110010010",
"011010011111001010000110",
"011010011110000101111110",
"011010011101000001111010",
"011010011011111101111010",
"011010011010111001111110",
"011010011001110110000111",
"011010011000110010010011",
"011010010111101110100100",
"011010010110101010111000",
"011010010101100111010001",
"011010010100100011101110",
"011010010011100000001111",
"011010010010011100110011",
"011010010001011001011100",
"011010010000010110001001",
"011010001111010010111010",
"011010001110001111101111",
"011010001101001100101000",
"011010001100001001100101",
"011010001011000110100110",
"011010001010000011101011",
"011010001001000000110101",
"011010000111111110000010",
"011010000110111011010011",
"011010000101111000101000",
"011010000100110110000001",
"011010000011110011011110",
"011010000010110000111111",
"011010000001101110100100",
"011010000000101100001101",
"011001111111101001111010",
"011001111110100111101011",
"011001111101100101100000",
"011001111100100011011001",
"011001111011100001010101",
"011001111010011111010110",
"011001111001011101011011",
"011001111000011011100011",
"011001110111011001110000",
"011001110110011000000000",
"011001110101010110010100",
"011001110100010100101101",
"011001110011010011001001",
"011001110010010001101001",
"011001110001010000001101",
"011001110000001110110101",
"011001101111001101100000",
"011001101110001100010000",
"011001101101001011000011",
"011001101100001001111011",
"011001101011001000110110",
"011001101010000111110101",
"011001101001000110111000",
"011001101000000101111111",
"011001100111000101001001",
"011001100110000100011000",
"011001100101000011101010",
"011001100100000011000000",
"011001100011000010011010",
"011001100010000001111000",
"011001100001000001011010",
"011001100000000000111111",
"011001011111000000101000",
"011001011110000000010110",
"011001011101000000000110",
"011001011011111111111011",
"011001011010111111110011",
"011001011001111111110000",
"011001011000111111110000",
"011001010111111111110100",
"011001010110111111111011",
"011001010110000000000110",
"011001010101000000010101",
"011001010100000000101000",
"011001010011000000111111",
"011001010010000001011001",
"011001010001000001110111",
"011001010000000010011001",
"011001001111000010111111",
"011001001110000011101000",
"011001001101000100010101",
"011001001100000101000110",
"011001001011000101111010",
"011001001010000110110011",
"011001001001000111101110",
"011001001000001000101110",
"011001000111001001110001",
"011001000110001010111000",
"011001000101001100000011",
"011001000100001101010001",
"011001000011001110100011",
"011001000010001111111001",
"011001000001010001010011",
"011001000000010010110000",
"011000111111010100010000",
"011000111110010101110101",
"011000111101010111011101",
"011000111100011001001001",
"011000111011011010111000",
"011000111010011100101011",
"011000111001011110100001",
"011000111000100000011100",
"011000110111100010011010",
"011000110110100100011011",
"011000110101100110100000",
"011000110100101000101001",
"011000110011101010110101",
"011000110010101101000101",
"011000110001101111011001",
"011000110000110001110000",
"011000101111110100001011",
"011000101110110110101001",
"011000101101111001001011",
"011000101100111011110000",
"011000101011111110011010",
"011000101011000001000110",
"011000101010000011110110",
"011000101001000110101010",
"011000101000001001100001",
"011000100111001100011100",
"011000100110001111011011",
"011000100101010010011101",
"011000100100010101100010",
"011000100011011000101011",
"011000100010011011111000",
"011000100001011111001000",
"011000100000100010011100",
"011000011111100101110011",
"011000011110101001001110",
"011000011101101100101100",
"011000011100110000001101",
"011000011011110011110011",
"011000011010110111011011",
"011000011001111011000111",
"011000011000111110110111",
"011000011000000010101010",
"011000010111000110100001",
"011000010110001010011011",
"011000010101001110011001",
"011000010100010010011010",
"011000010011010110011110",
"011000010010011010100110",
"011000010001011110110010",
"011000010000100011000001",
"011000001111100111010011",
"011000001110101011101001",
"011000001101110000000010",
"011000001100110100011111",
"011000001011111000111111",
"011000001010111101100010",
"011000001010000010001001",
"011000001001000110110100",
"011000001000001011100001",
"011000000111010000010011",
"011000000110010101000111",
"011000000101011001111111",
"011000000100011110111011",
"011000000011100011111001",
"011000000010101000111100",
"011000000001101110000001",
"011000000000110011001010",
"010111111111111000010110",
"010111111110111101100110",
"010111111110000010111001",
"010111111101001000010000",
"010111111100001101101001",
"010111111011010011000111",
"010111111010011000100111",
"010111111001011110001011",
"010111111000100011110010",
"010111110111101001011101",
"010111110110101111001011",
"010111110101110100111100",
"010111110100111010110000",
"010111110100000000101000",
"010111110011000110100100",
"010111110010001100100010",
"010111110001010010100100",
"010111110000011000101001",
"010111101111011110110010",
"010111101110100100111101",
"010111101101101011001100",
"010111101100110001011111",
"010111101011110111110100",
"010111101010111110001101",
"010111101010000100101010",
"010111101001001011001001",
"010111101000010001101100",
"010111100111011000010010",
"010111100110011110111011",
"010111100101100101101000",
"010111100100101100011000",
"010111100011110011001011",
"010111100010111010000001",
"010111100010000000111011",
"010111100001000111111000",
"010111100000001110111000",
"010111011111010101111011",
"010111011110011101000001",
"010111011101100100001011",
"010111011100101011011000",
"010111011011110010101000",
"010111011010111001111100",
"010111011010000001010011",
"010111011001001000101100",
"010111011000010000001010",
"010111010111010111101010",
"010111010110011111001101",
"010111010101100110110100",
"010111010100101110011110",
"010111010011110110001011",
"010111010010111101111011",
"010111010010000101101110",
"010111010001001101100101",
"010111010000010101011111",
"010111001111011101011100",
"010111001110100101011100",
"010111001101101101011111",
"010111001100110101100110",
"010111001011111101101111",
"010111001011000101111100",
"010111001010001110001100",
"010111001001010110011111",
"010111001000011110110101",
"010111000111100111001110",
"010111000110101111101011",
"010111000101111000001010",
"010111000101000000101101",
"010111000100001001010011",
"010111000011010001111011",
"010111000010011010100111",
"010111000001100011010111",
"010111000000101100001001",
"010110111111110100111110",
"010110111110111101110111",
"010110111110000110110010",
"010110111101001111110001",
"010110111100011000110010",
"010110111011100001110111",
"010110111010101010111111",
"010110111001110100001010",
"010110111000111101011000",
"010110111000000110101001",
"010110110111001111111101",
"010110110110011001010101",
"010110110101100010101111",
"010110110100101100001100",
"010110110011110101101101",
"010110110010111111010000",
"010110110010001000110111",
"010110110001010010100000",
"010110110000011100001101",
"010110101111100101111100",
"010110101110101111101111",
"010110101101111001100101",
"010110101101000011011101",
"010110101100001101011001",
"010110101011010111011000",
"010110101010100001011001",
"010110101001101011011110",
"010110101000110101100110",
"010110100111111111110001",
"010110100111001001111110",
"010110100110010100001111",
"010110100101011110100011",
"010110100100101000111010",
"010110100011110011010011",
"010110100010111101110000",
"010110100010001000010000",
"010110100001010010110010",
"010110100000011101011000",
"010110011111101000000001",
"010110011110110010101100",
"010110011101111101011011",
"010110011101001000001100",
"010110011100010011000001",
"010110011011011101111000",
"010110011010101000110010",
"010110011001110011110000",
"010110011000111110110000",
"010110011000001001110011",
"010110010111010100111001",
"010110010110100000000010",
"010110010101101011001110",
"010110010100110110011101",
"010110010100000001101111",
"010110010011001101000011",
"010110010010011000011011",
"010110010001100011110101",
"010110010000101111010011",
"010110001111111010110011",
"010110001111000110010110",
"010110001110010001111101",
"010110001101011101100110",
"010110001100101001010010",
"010110001011110101000000",
"010110001011000000110010",
"010110001010001100100111",
"010110001001011000011110",
"010110001000100100011000",
"010110000111110000010110",
"010110000110111100010110",
"010110000110001000011001",
"010110000101010100011110",
"010110000100100000100111",
"010110000011101100110010",
"010110000010111001000001",
"010110000010000101010010",
"010110000001010001100110",
"010110000000011101111101",
"010101111111101010010111",
"010101111110110110110011",
"010101111110000011010011",
"010101111101001111110101",
"010101111100011100011010",
"010101111011101001000010",
"010101111010110101101100",
"010101111010000010011010",
"010101111001001111001010",
"010101111000011011111101",
"010101110111101000110011",
"010101110110110101101100",
"010101110110000010100111",
"010101110101001111100110",
"010101110100011100100111",
"010101110011101001101011",
"010101110010110110110001",
"010101110010000011111011",
"010101110001010001000111",
"010101110000011110010110",
"010101101111101011101000",
"010101101110111000111101",
"010101101110000110010100",
"010101101101010011101110",
"010101101100100001001011",
"010101101011101110101011",
"010101101010111100001101",
"010101101010001001110010",
"010101101001010111011010",
"010101101000100101000101",
"010101100111110010110010",
"010101100111000000100010",
"010101100110001110010101",
"010101100101011100001010",
"010101100100101010000011",
"010101100011110111111110",
"010101100011000101111011",
"010101100010010011111100",
"010101100001100001111111",
"010101100000110000000101",
"010101011111111110001110",
"010101011111001100011001",
"010101011110011010100111",
"010101011101101000111000",
"010101011100110111001011",
"010101011100000101100001",
"010101011011010011111010",
"010101011010100010010110",
"010101011001110000110100",
"010101011000111111010101",
"010101011000001101111000",
"010101010111011100011111",
"010101010110101011000111",
"010101010101111001110011",
"010101010101001000100001",
"010101010100010111010010",
"010101010011100110000110",
"010101010010110100111100",
"010101010010000011110101",
"010101010001010010110001",
"010101010000100001101111",
"010101001111110000110000",
"010101001110111111110011",
"010101001110001110111001",
"010101001101011110000010",
"010101001100101101001101",
"010101001011111100011011",
"010101001011001011101100",
"010101001010011010111111",
"010101001001101010010101",
"010101001000111001101110",
"010101001000001001001001",
"010101000111011000100111",
"010101000110101000000111",
"010101000101110111101010",
"010101000101000111010000",
"010101000100010110111000",
"010101000011100110100011",
"010101000010110110010000",
"010101000010000110000000",
"010101000001010101110011",
"010101000000100101101000",
"010100111111110101100000",
"010100111111000101011010",
"010100111110010101010111",
"010100111101100101010111",
"010100111100110101011001",
"010100111100000101011110",
"010100111011010101100101",
"010100111010100101101111",
"010100111001110101111011",
"010100111001000110001010",
"010100111000010110011011",
"010100110111100110101111",
"010100110110110111000110",
"010100110110000111011111",
"010100110101010111111011",
"010100110100101000011001",
"010100110011111000111010",
"010100110011001001011101",
"010100110010011010000011",
"010100110001101010101011",
"010100110000111011010110",
"010100110000001100000100",
"010100101111011100110100",
"010100101110101101100110",
"010100101101111110011011",
"010100101101001111010011",
"010100101100100000001101",
"010100101011110001001001",
"010100101011000010001000",
"010100101010010011001010",
"010100101001100100001110",
"010100101000110101010100",
"010100101000000110011101",
"010100100111010111101001",
"010100100110101000110111",
"010100100101111010000111",
"010100100101001011011010",
"010100100100011100110000",
"010100100011101110001000",
"010100100010111111100010",
"010100100010010000111111",
"010100100001100010011111",
"010100100000110100000000",
"010100100000000101100101",
"010100011111010111001011",
"010100011110101000110101",
"010100011101111010100000",
"010100011101001100001110",
"010100011100011101111111",
"010100011011101111110010",
"010100011011000001101000",
"010100011010010011100000",
"010100011001100101011010",
"010100011000110111010111",
"010100011000001001010110",
"010100010111011011011000",
"010100010110101101011100",
"010100010101111111100010",
"010100010101010001101011",
"010100010100100011110111",
"010100010011110110000100",
"010100010011001000010101",
"010100010010011010100111",
"010100010001101100111100",
"010100010000111111010100",
"010100010000010001101110",
"010100001111100100001010",
"010100001110110110101001",
"010100001110001001001010",
"010100001101011011101101",
"010100001100101110010011",
"010100001100000000111011",
"010100001011010011100110",
"010100001010100110010011",
"010100001001111001000010",
"010100001001001011110100",
"010100001000011110101000",
"010100000111110001011111",
"010100000111000100011000",
"010100000110010111010011",
"010100000101101010010001",
"010100000100111101010001",
"010100000100010000010011",
"010100000011100011011000",
"010100000010110110011111",
"010100000010001001101000",
"010100000001011100110100",
"010100000000110000000010",
"010100000000000011010011",
"010011111111010110100101",
"010011111110101001111011",
"010011111101111101010010",
"010011111101010000101100",
"010011111100100100001000",
"010011111011110111100111",
"010011111011001011001000",
"010011111010011110101011",
"010011111001110010010000",
"010011111001000101111000",
"010011111000011001100010",
"010011110111101101001111",
"010011110111000000111101",
"010011110110010100101110",
"010011110101101000100010",
"010011110100111100011000",
"010011110100010000001111",
"010011110011100100001010",
"010011110010111000000110",
"010011110010001100000101",
"010011110001100000000110",
"010011110000110100001010",
"010011110000001000010000",
"010011101111011100011000",
"010011101110110000100010",
"010011101110000100101111",
"010011101101011000111110",
"010011101100101101001111",
"010011101100000001100010",
"010011101011010101111000",
"010011101010101010010000",
"010011101001111110101010",
"010011101001010011000111",
"010011101000100111100101",
"010011100111111100000110",
"010011100111010000101010",
"010011100110100101001111",
"010011100101111001110111",
"010011100101001110100001",
"010011100100100011001101",
"010011100011110111111100",
"010011100011001100101101",
"010011100010100001100000",
"010011100001110110010101",
"010011100001001011001100",
"010011100000100000000110",
"010011011111110101000010",
"010011011111001010000000",
"010011011110011111000001",
"010011011101110100000011",
"010011011101001001001000",
"010011011100011110001111",
"010011011011110011011000",
"010011011011001000100100",
"010011011010011101110010",
"010011011001110011000001",
"010011011001001000010100",
"010011011000011101101000",
"010011010111110010111110",
"010011010111001000010111",
"010011010110011101110010",
"010011010101110011001111",
"010011010101001000101110",
"010011010100011110010000",
"010011010011110011110100",
"010011010011001001011001",
"010011010010011111000001",
"010011010001110100101100",
"010011010001001010011000",
"010011010000100000000111",
"010011001111110101110111",
"010011001111001011101010",
"010011001110100001011111",
"010011001101110111010111",
"010011001101001101010000",
"010011001100100011001100",
"010011001011111001001001",
"010011001011001111001001",
"010011001010100101001011",
"010011001001111011001111",
"010011001001010001010110",
"010011001000100111011110",
"010011000111111101101001",
"010011000111010011110110",
"010011000110101010000101",
"010011000110000000010110",
"010011000101010110101001",
"010011000100101100111110",
"010011000100000011010110",
"010011000011011001101111",
"010011000010110000001011",
"010011000010000110101001",
"010011000001011101001001",
"010011000000110011101011",
"010011000000001010001111",
"010010111111100000110110",
"010010111110110111011110",
"010010111110001110001000",
"010010111101100100110101",
"010010111100111011100100",
"010010111100010010010101",
"010010111011101001001000",
"010010111010111111111101",
"010010111010010110110100",
"010010111001101101101101",
"010010111001000100101001",
"010010111000011011100110",
"010010110111110010100110",
"010010110111001001100111",
"010010110110100000101011",
"010010110101110111110001",
"010010110101001110111001",
"010010110100100110000011",
"010010110011111101001111",
"010010110011010100011101",
"010010110010101011101101",
"010010110010000010111111",
"010010110001011010010011",
"010010110000110001101010",
"010010110000001001000010",
"010010101111100000011101",
"010010101110110111111001",
"010010101110001111011000",
"010010101101100110111001",
"010010101100111110011011",
"010010101100010110000000",
"010010101011101101100111",
"010010101011000101010000",
"010010101010011100111011",
"010010101001110100101000",
"010010101001001100010110",
"010010101000100100001000",
"010010100111111011111011",
"010010100111010011110000",
"010010100110101011100111",
"010010100110000011100000",
"010010100101011011011011",
"010010100100110011011000",
"010010100100001011010111",
"010010100011100011011001",
"010010100010111011011100",
"010010100010010011100001",
"010010100001101011101000",
"010010100001000011110010",
"010010100000011011111101",
"010010011111110100001010",
"010010011111001100011010",
"010010011110100100101011",
"010010011101111100111110",
"010010011101010101010100",
"010010011100101101101011",
"010010011100000110000100",
"010010011011011110100000",
"010010011010110110111101",
"010010011010001111011100",
"010010011001100111111101",
"010010011001000000100001",
"010010011000011001000110",
"010010010111110001101101",
"010010010111001010010110",
"010010010110100011000001",
"010010010101111011101110",
"010010010101010100011110",
"010010010100101101001111",
"010010010100000110000010",
"010010010011011110110111",
"010010010010110111101110",
"010010010010010000100111",
"010010010001101001100001",
"010010010001000010011110",
"010010010000011011011101",
"010010001111110100011110",
"010010001111001101100001",
"010010001110100110100101",
"010010001101111111101100",
"010010001101011000110100",
"010010001100110001111111",
"010010001100001011001011",
"010010001011100100011010",
"010010001010111101101010",
"010010001010010110111100",
"010010001001110000010000",
"010010001001001001100110",
"010010001000100010111111",
"010010000111111100011000",
"010010000111010101110100",
"010010000110101111010010",
"010010000110001000110010",
"010010000101100010010100",
"010010000100111011110111",
"010010000100010101011101",
"010010000011101111000100",
"010010000011001000101101",
"010010000010100010011000",
"010010000001111100000110",
"010010000001010101110101",
"010010000000101111100101",
"010010000000001001011000",
"010001111111100011001101",
"010001111110111101000100",
"010001111110010110111100",
"010001111101110000110111",
"010001111101001010110011",
"010001111100100100110001",
"010001111011111110110001",
"010001111011011000110011",
"010001111010110010110111",
"010001111010001100111101",
"010001111001100111000100",
"010001111001000001001110",
"010001111000011011011001",
"010001110111110101100110",
"010001110111001111110101",
"010001110110101010000110",
"010001110110000100011001",
"010001110101011110101110",
"010001110100111001000101",
"010001110100010011011101",
"010001110011101101110111",
"010001110011001000010011",
"010001110010100010110001",
"010001110001111101010001",
"010001110001010111110011",
"010001110000110010010111",
"010001110000001100111100",
"010001101111100111100011",
"010001101111000010001100",
"010001101110011100110111",
"010001101101110111100100",
"010001101101010010010011",
"010001101100101101000011",
"010001101100000111110101",
"010001101011100010101010",
"010001101010111101011111",
"010001101010011000010111",
"010001101001110011010001",
"010001101001001110001100",
"010001101000101001001010",
"010001101000000100001001",
"010001100111011111001010",
"010001100110111010001100",
"010001100110010101010001",
"010001100101110000010111",
"010001100101001011011111",
"010001100100100110101001",
"010001100100000001110101",
"010001100011011101000011",
"010001100010111000010010",
"010001100010010011100011",
"010001100001101110110110",
"010001100001001010001011",
"010001100000100101100010",
"010001100000000000111010",
"010001011111011100010101",
"010001011110110111110001",
"010001011110010011001110",
"010001011101101110101110",
"010001011101001010001111",
"010001011100100101110010",
"010001011100000001010111",
"010001011011011100111110",
"010001011010111000100111",
"010001011010010100010001",
"010001011001101111111101",
"010001011001001011101011",
"010001011000100111011010",
"010001011000000011001100",
"010001010111011110111111",
"010001010110111010110100",
"010001010110010110101010",
"010001010101110010100011",
"010001010101001110011101",
"010001010100101010011001",
"010001010100000110010111",
"010001010011100010010110",
"010001010010111110010111",
"010001010010011010011010",
"010001010001110110011111",
"010001010001010010100110",
"010001010000101110101110",
"010001010000001010111000",
"010001001111100111000011",
"010001001111000011010001",
"010001001110011111100000",
"010001001101111011110001",
"010001001101011000000100",
"010001001100110100011000",
"010001001100010000101110",
"010001001011101101000110",
"010001001011001001100000",
"010001001010100101111011",
"010001001010000010011000",
"010001001001011110110111",
"010001001000111011010111",
"010001001000010111111010",
"010001000111110100011110",
"010001000111010001000011",
"010001000110101101101011",
"010001000110001010010100",
"010001000101100110111110",
"010001000101000011101011",
"010001000100100000011001",
"010001000011111101001001",
"010001000011011001111011",
"010001000010110110101110",
"010001000010010011100011",
"010001000001110000011010",
"010001000001001101010010",
"010001000000101010001101",
"010001000000000111001000",
"010000111111100100000110",
"010000111111000001000101",
"010000111110011110000110",
"010000111101111011001001",
"010000111101011000001101",
"010000111100110101010011",
"010000111100010010011011",
"010000111011101111100100",
"010000111011001100101111",
"010000111010101001111100",
"010000111010000111001010",
"010000111001100100011010",
"010000111001000001101100",
"010000111000011110111111",
"010000110111111100010100",
"010000110111011001101011",
"010000110110110111000011",
"010000110110010100011101",
"010000110101110001111001",
"010000110101001111010111",
"010000110100101100110110",
"010000110100001010010110",
"010000110011100111111001",
"010000110011000101011101",
"010000110010100011000010",
"010000110010000000101010",
"010000110001011110010011",
"010000110000111011111101",
"010000110000011001101010",
"010000101111110111011000",
"010000101111010101000111",
"010000101110110010111000",
"010000101110010000101011",
"010000101101101110100000",
"010000101101001100010110",
"010000101100101010001101",
"010000101100001000000111",
"010000101011100110000010",
"010000101011000011111111",
"010000101010100001111101",
"010000101001111111111101",
"010000101001011101111110",
"010000101000111100000001",
"010000101000011010000110",
"010000100111111000001101",
"010000100111010110010101",
"010000100110110100011110",
"010000100110010010101001",
"010000100101110000110110",
"010000100101001111000101",
"010000100100101101010101",
"010000100100001011100111",
"010000100011101001111010",
"010000100011001000001111",
"010000100010100110100101",
"010000100010000100111101",
"010000100001100011010111",
"010000100001000001110011",
"010000100000100000001111",
"010000011111111110101110",
"010000011111011101001110",
"010000011110111011110000",
"010000011110011010010011",
"010000011101111000111000",
"010000011101010111011110",
"010000011100110110000110",
"010000011100010100110000",
"010000011011110011011011",
"010000011011010010001000",
"010000011010110000110111",
"010000011010001111100111",
"010000011001101110011000",
"010000011001001101001011",
"010000011000101100000000",
"010000011000001010110110",
"010000010111101001101110",
"010000010111001000101000",
"010000010110100111100010",
"010000010110000110011111",
"010000010101100101011101",
"010000010101000100011101",
"010000010100100011011110",
"010000010100000010100001",
"010000010011100001100101",
"010000010011000000101011",
"010000010010011111110011",
"010000010001111110111100",
"010000010001011110000110",
"010000010000111101010010",
"010000010000011100100000",
"010000001111111011101111",
"010000001111011011000000",
"010000001110111010010011",
"010000001110011001100110",
"010000001101111000111100",
"010000001101011000010011",
"010000001100110111101011",
"010000001100010111000101",
"010000001011110110100001",
"010000001011010101111110",
"010000001010110101011101",
"010000001010010100111101",
"010000001001110100011111",
"010000001001010100000010",
"010000001000110011100111",
"010000001000010011001101",
"010000000111110010110101",
"010000000111010010011110",
"010000000110110010001001",
"010000000110010001110101",
"010000000101110001100011",
"010000000101010001010010",
"010000000100110001000011",
"010000000100010000110110",
"010000000011110000101010",
"010000000011010000011111",
"010000000010110000010110",
"010000000010010000001111",
"010000000001110000001001",
"010000000001010000000100",
"010000000000110000000001",
"010000000000010000000000"
);

end package fp_inv_table;
