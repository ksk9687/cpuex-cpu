-- @module : cpu_top
-- @author : ksk
-- @date   : 2009/10/06


library ieee;
use ieee.std_logic_1164.all;

entity cpu_top is 
port (
    clk			: in	  std_logic
    
    
    ); 
     
end cpu_top;     
        

architecture synth of cpu_top is
               
begin  

end synth;








