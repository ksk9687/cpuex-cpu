--�@������

-- @module : mem
-- @author : ksk
-- @date   : 2009/10/06



library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library work;
use work.instruction.all;

entity mem is 
port (
    clk,sramcclk,sramclk	: in	  std_logic;
    
    pc : in std_logic_vector(31 downto 0);
    ls_address : in std_logic_vector(31 downto 0);
    load_store : in std_logic_vector(1 downto 0);
    write_data : in std_logic_vector(31 downto 0);
    read_inst,read_data : out std_logic_vector(31 downto 0);
    read_data_ready : out std_logic
    
    
	--SRAM
	;SRAMAA : out  STD_LOGIC_VECTOR (19 downto 0)	--�A�h���X
	;SRAMIOA : inout  STD_LOGIC_VECTOR (31 downto 0)	--�f�[�^
	;SRAMIOPA : inout  STD_LOGIC_VECTOR (3 downto 0) --�p���e�B�[
	
	;SRAMRWA : out  STD_LOGIC	--read=>1,write=>0
	;SRAMBWA : out  STD_LOGIC_VECTOR (3 downto 0)--�������݃o�C�g�̎w��

	;SRAMCLKMA0 : out  STD_LOGIC	--SRAM�N���b�N
	;SRAMCLKMA1 : out  STD_LOGIC	--SRAM�N���b�N
	
	;SRAMADVLDA : out  STD_LOGIC	--�o�[�X�g�A�N�Z�X
	;SRAMCEA : out  STD_LOGIC --clock enable
	
	;SRAMCELA1X : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���
	;SRAMCEHA1X : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���
	;SRAMCEA2X : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���
	;SRAMCEA2 : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���

	;SRAMLBOA : out  STD_LOGIC	--�o�[�X�g�A�N�Z�X��
	;SRAMXOEA : out  STD_LOGIC	--IO�o�̓C�l�[�u��
	;SRAMZZA : out  STD_LOGIC	--�X���[�v���[�h�ɓ���
    ); 
     
     constant sleep : std_logic_vector(31 downto 0):= op_halt&"00"&"00000000"&"00000000"&"00000000";
end mem;
        

architecture synth of mem is
	type mem_state is (init,
	inst,inst_w1,inst_w2,inst_w3,inst_w4,data,
	data_w1,data_w2,data_w3,data_w4,load_end
	);
	signal state : mem_state := init;
	signal count : std_logic_vector(31 downto 0) := (others => '0');
	
	signal RW : std_logic := '0';
	signal DATAIN : std_logic_vector(31 downto 0) := (others => '0');
	signal DATAOUT : std_logic_vector(31 downto 0) := (others => '0');
	signal ADDR : std_logic_vector(19 downto 0) := (others => '0');
	
    type ram_type is array (0 to 15) of std_logic_vector (31 downto 0); 
	signal RAM : ram_type :=
--	(--fib10
--	op_li & "00000" & "00000" & x"0000",
--	op_li & "00000" & "00001" & x"0000",
--	op_li & "00000" & "00010" & x"0001",
--	op_li & "00000" & "00011" & x"000A",
--	
--	op_li & "00000" & "00100" & x"0001",
--	op_add & "00001" & "00010" & "00000" & "00000000000",
--	op_addi & "00010" & "00001" & x"0000",
--	op_addi & "00000" & "00010" & x"0000",
--	
--	op_addi & "00011" & "00011" & x"FFFF",
--	op_cmp & "00011" & "00100" & "00101" & "00000000000",
--	op_jmp & "00101" & "00011" & x"FFFB",-- -5\
--	--op_write & "00000" & "00000" & x"0000",
--	op_store & "00011" & "00000" & x"0000",
--
--
--	--op_store & "00011" & "00000" & x"0001",
--	--op_nop & "00000" & "00000" & x"0000",
--	op_load & "00011" & "00000" & x"0000",
--	op_write & "00000" & "00000" & x"0000",
--	--op_halt & "00000" & "00000" & x"0000",
--	--op_halt & "00000" & "00000" & x"0000",
--	op_halt & "00000" & "00000" & x"0000",
--	op_halt & "00000" & "00000" & x"0000"
--	);
		(--ls
	op_li & "00000" & "00000" & op_li & "00000" & "00000",
	op_sll & "00000" & "00000" & x"0010",
	op_addi & "00000" & "00000" & x"0033",
	op_li & "00000" & "00001" & x"0000",
	
	op_li & "00000" & "00010" & x"0007",
	op_load & "00001" & "00010" & x"0008",
	op_write & "00010" & "00000" & x"0000",
	op_halt & "00000" & "00000" & x"0000",
	
	op_halt & "00000" & "00000" & x"00"&"00011001",
	op_halt & "00000" & "00000" & x"0000",
	op_halt & "00000" & "00000" & x"0000",
	op_halt & "00000" & "00000" & x"0000",
	
	op_halt & "00000" & "00000" & x"0000",
	op_halt & "00000" & "00000" & x"0000",
	op_halt & "00000" & "00000" & x"0000",
	op_halt & "00000" & "00000" & x"0000"
	);
	component sram_controller is
    Port (
		CLK : in STD_LOGIC
		;SRAMCLK : in STD_LOGIC
		;ADDR    : in  std_logic_vector(19 downto 0)
		;DATAIN  : in  std_logic_vector(31 downto 0)
		;DATAOUT : out std_logic_vector(31 downto 0)
		;RW      : in  std_logic
		--SRAM
		;SRAMAA : out  STD_LOGIC_VECTOR (19 downto 0)	--�A�h���X
		;SRAMIOA : inout  STD_LOGIC_VECTOR (31 downto 0)	--�f�[�^
		;SRAMIOPA : inout  STD_LOGIC_VECTOR (3 downto 0) --�p���e�B�[
		
		;SRAMRWA : out  STD_LOGIC	--read=>1,write=>0
		;SRAMBWA : out  STD_LOGIC_VECTOR (3 downto 0)--�������݃o�C�g�̎w��

		;SRAMCLKMA0 : out  STD_LOGIC	--SRAM�N���b�N
		;SRAMCLKMA1 : out  STD_LOGIC	--SRAM�N���b�N
		
		;SRAMADVLDA : out  STD_LOGIC	--�o�[�X�g�A�N�Z�X
		;SRAMCEA : out  STD_LOGIC --clock enable
		
		;SRAMCELA1X : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���
		;SRAMCEHA1X : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���
		;SRAMCEA2X : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���
		;SRAMCEA2 : out  STD_LOGIC	--SRAM�𓮍삳���邩�ǂ���
		
		;SRAMLBOA : out  STD_LOGIC	--�o�[�X�g�A�N�Z�X��
		;SRAMXOEA : out  STD_LOGIC	--IO�o�̓C�l�[�u��
		;SRAMZZA : out  STD_LOGIC	--�X���[�v���[�h�ɓ���
	);
	end component;
begin

	--�Ƃ肠�������URAM���������Ƃ��ė��p����
	  
--	--�f�[�^
--	process (clk)
--	begin
--	    if rising_edge(clk) then
--	        if load_store = '1' then
--	            RAM(conv_integer(ls_address(3 downto 0))) <= write_data;
--	        end if;
--	    end if;
--	end process;
--	read_data <= RAM(conv_integer(ls_address(3 downto 0)));
--	
--	-- ����
--	read_inst <= RAM(conv_integer(pc(3 downto 0)));


	
	ADDR <= count(19 downto 0) when state = init else
	pc(19 downto 0) when state = inst else
	ls_address(19 downto 0) when state = data else
	(others => '0');
	
	DATAIN <= RAM(conv_integer(count(3 downto 0))) when state = init else
	write_data when (state = data) else
	(others => '0');
	
	RW <= '0' when state = init else--w
	(not load_store(0)) when state = data else
	'1';
	
	read_inst <= DATAOUT when state = data else
	sleep;
	
	read_data_ready <= '1' when state = load_end else
	'0';
	
	read_data <= DATAOUT when state = inst else
	"010101010101"&"0101010101"&"0101010101";
	
	
	process(clk)
	begin
	if rising_edge(clk) then
		if state = init then
			if count(4 downto 0) = "10000" then
				state <= inst;
			else
				state <= state;
			end if;
		elsif state = inst then 
			state <= inst_w1;
		elsif state = inst_w1 then 
			state <= inst_w2;
		elsif state = inst_w2 then 
			state <= inst_w3;
		elsif state = inst_w3 then 
			state <= data;
		elsif state = inst_w4 then
			state <= data;
		elsif state = data then
			if (load_store = "10") then--Load�����L�т�
				state <= data_w1;
			else
				state <= inst;
			end if;
		elsif state = data_w1 then
			state <= data_w2;
		elsif state = data_w2 then
			state <= data_w3;
		elsif state = data_w3 then
			state <= inst;
		elsif state = load_end then
			state <= inst;
		end if;
		count <= count + '1';
	end if;
	end process;

	SRAMC : sram_controller port map(
		 sramcclk
		,sramclk
		,ADDR
		,DATAIN
		,DATAOUT
		,RW
		,SRAMAA,SRAMIOA,SRAMIOPA
		,SRAMRWA,SRAMBWA
		,SRAMCLKMA0,SRAMCLKMA1
		,SRAMADVLDA,SRAMCEA
		,SRAMCELA1X,SRAMCEHA1X,SRAMCEA2X,SRAMCEA2
		,SRAMLBOA,SRAMXOEA,SRAMZZA
	);

end synth;








