library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;

library unisim;
use unisim.vcomponents.all;

entity FP_ADD_TESTER is
  port (
    clkin  : in  std_logic;
    ledout : out std_logic_vector(1 downto 0));
end FP_ADD_TESTER;


architecture STRUCTURE of FP_ADD_TESTER is

  component FP_ADD
    port (
      A, B : in  std_logic_vector(31 downto 0); 
      O    : out std_logic_vector(31 downto 0));
  end component;



  constant n : integer := 100;
  subtype float is std_logic_vector(31 downto 0);
  type table is array(0 to n-1) of float;

  constant table_a : table := (
    "00000000000000000000000000000000",
    "11010111010111111000100101000101",
    "00100001011100010110000111000100",
    "00110100101101111001010100100111",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "01110100011101110110101101011001",
    "11101100101000100011100000000000",
    "11101000000001000011100111110111",
    "00001100011011111111000111000010",
    "10010010001001001100011110101101",
    "00111011111001110010101010001010",
    "00100010111010100010101011111001",
    "01101000001100101100111010101000",
    "01001111010001110111100010010100",
    "01111011110111100010010101001110",
    "01011100000100011010101110101001",
    "00011100000001101111000011111110",
    "01100010011000011011101110111001",
    "00100111100110001010101111011000",
    "00111001010100011110111110011111",
    "01101101000000010100111111001011",
    "01110010101001100000010010111100",
    "10111011000101100001101111011101",
    "00000110000000100110100100010011",
    "10111000101111010010001110000100",
    "10111001111001011000000000100011",
    "01001110001011011111111111001001",
    "10110011011010100110110100100111",
    "01011101001011111111001101001011",
    "10101110010010110100000101010011",
    "00100011010100101000110111000110",
    "00111011101111000001000011000000",
    "10010100011111000100000101001100",
    "11000001011001110001111000101000",
    "10001111000110001001110011010111",
    "10000011011101110100001000111101",
    "11011110000001100010010111011100",
    "10111010000011111011001010111100",
    "11111101101100111010000110100001",
    "01011010011011100101110110111010",
    "01110000010001111011100001110100",
    "11000101101010000011100111100000",
    "11101100010000001100110010111100",
    "10100010100010110000001101001110",
    "10110110010010111101111110000011",
    "10001110100000100011000100001101",
    "10101100011000110000011111000010",
    "11010010110101010001011101111011",
    "10100000011011000001101010011010",
    "11100100110101011100001101101101",
    "10110000111000100100110100011111",
    "01000111011011110111111010111100",
    "01001111100100100001110101110101",
    "10101011111111110000010001000001",
    "10100001111101010101110101101011",
    "11111100110010010101010111101011",
    "00110011000000111001110011100011",
    "00010101111011000001010111000001",
    "01110100010110000010001111000110",
    "01001101110100100010000111101111",
    "01110010111110001000000110001000",
    "00110011001011000111011000111010",
    "00111100101101100011000110000001",
    "10111001110111101011000111010101",
    "11101110010111001100111100001011",
    "10111000001101101101001000010001",
    "10110001110000101001100000010010",
    "00001111100001100011011101100101",
    "10000001101110101111000100011111",
    "00011111001110111110010111100110",
    "00001001101110000000111100010001",
    "11111010000111100110101011000010",
    "01100010100100111100101001111110",
    "00001111010101010011000011111010",
    "01110011001100001100001011001000",
    "11011011110011010110011010100011",
    "10110011101100101101010010111001",
    "11001111010010000111010010011101",
    "10110100101011110101111010010110",
    "10011110101100110100101101000011",
    "01111001010010001101101010001000",
    "00011010010100000100001001000111",
    "10100100010101011110010100100000",
    "10000011110111111001111100001111",
    "11100000010110100101100011110110",
    "10100010010110010010011010011010",
    "01111101010001011010111100011010",
    "01111000001010011101010010100110",
    "01101110100010100101111010000011",
    "01011011000001010101010001101110",
    "11110011010000010111100000101000",
    "10110010110001000101011011000001",
    "01011011110100101101001000110101",
    "00010011110010010000111110110001",
    "01001001010010011011100000010111",
    "10110011110010001111101100010101",
    "01110101110000100110011100011010",
    "10110001011010110111110010110001");

  constant table_b : table := (
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "01111001100000000001100111010011",
    "11001000011010010001110110111110",
    "11011000100111000100011000001010",
    "11110100011101110110101101011001",
    "01101100101000100011100000000000",
    "01101000000001000011100111110111",
    "10001100011011111111000111000010",
    "00010010001001001100011110101101",
    "10111011111001110010101010001010",
    "10100010111010100010101011111001",
    "11101000001100101100111010101000",
    "11001111010001110111100010010100",
    "11111011110111100010010101001110",
    "10100110111000110101010010001010",
    "01011101011011001111100001101010",
    "01001101010110110011000000011010",
    "10000110101010010011111111001001",
    "10000001001011001011011010000001",
    "10111111110011000110001000000110",
    "10010101110100011000111000001001",
    "10001111101101010010011001100100",
    "11011100111111001100010000110010",
    "11000001001111101100011100101011",
    "00001011100001110000110010100000",
    "10100010011101100111111011111101",
    "11000111011010101101100001111011",
    "01110100000110010101010000011001",
    "01001010000011101110110010110011",
    "00100001001101011011100001000001",
    "01000110000100101011110011100000",
    "01001100001101000100111000101111",
    "01001010001010111001000111011011",
    "01011101110010101101001010111000",
    "00110101000101010111010011000110",
    "11111001111100001100011011011110",
    "00011010110111010101101000110100",
    "11100110111000001011110110011101",
    "01010000110110101001001111010100",
    "01111110000111110100001101100010",
    "00111111100011000110101011001110",
    "01011011011100011001000111101110",
    "11000110101010101100111110011101",
    "10001001000001001111100110010101",
    "11111111010001110111011111100111",
    "11110110110000100001101111100100",
    "01001111111110001101010001110000",
    "10101011110101000011101111100011",
    "01010111101100110001101110011100",
    "10100010010101111011000010110000",
    "00101000110100011110010011100110",
    "11011100010011101001000000100011",
    "10100000010111101000000110000010",
    "10011001101101100100010000111010",
    "00001111000000110111001110000110",
    "01001100110000101011011011100110",
    "00110001000110100000100101111111",
    "01111110110001010001000000110011",
    "00111001001011001011010110011011",
    "00000101100111011001101010001011",
    "01010011000110100000011110110110",
    "10011000010001001110001111000000",
    "01100001011110100010011000010101",
    "10110100011000011011011100001011",
    "10111111101110011111001101011110",
    "10010100001010110110000010001111",
    "10001000100101000000111100001101",
    "01000011001111000000110101101001",
    "11010100010100100010100111110011",
    "01010010111110010000000000010010",
    "10011011110111110111100001010001",
    "00011110011001110001111100110010",
    "00010100100110101110011111110111",
    "11100011010110111011100100111110",
    "00001000101110010100100011111110",
    "10011001000010101100000001100110",
    "11011010000000010011110001000101",
    "01111010111001001000010100000010",
    "11010101100101010000001000010110",
    "01001100110110011100011111010001",
    "01000001001101011000011010101101",
    "11100001001000011100110101010100",
    "11010000110010100011011110100000",
    "00110111000000111100011110100010",
    "00001010010011011000011001001101",
    "10001000100100110000100010001101",
    "00011001011001001101010110101111",
    "00111110111110000000000110111111",
    "01001111111011010001011111110000",
    "01101000010000010110000001110001",
    "00101010101000110100111001101100",
    "00010111110111101011110100101001",
    "10011010011111111000100001011000",
    "11010101100101010100101000010010",
    "00010010001110100000010111111000",
    "10101011001001011111101101111101",
    "11011000001101101100101001000001");

  constant table_o : table := (
    "00000000000000000000000000000000",
    "11010111010111111000100101000101",
    "00100001011100010110000111000100",
    "00110100101101111001010100100111",
    "01111001100000000001100111010011",
    "11001000011010010001110110111110",
    "11011000100111000100011000001010",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "01011100000100011010101110101001",
    "01011101011011001111100001101010",
    "01100010011000011011101110111001",
    "00100111100110001010101111011000",
    "00111001010100011110111110011111",
    "01101101000000010100111111001011",
    "01110010101001100000010010111100",
    "10111011000101100001101111011101",
    "11011100111111001100010000110010",
    "11000001001111101100011110001001",
    "10111001111001011000000000100011",
    "01001110001011011111111111001001",
    "11000111011010101101100001111011",
    "01110100000110010101010000011001",
    "01001010000011101110110010110011",
    "00100011010111011110100101001010",
    "01000110000100101011110011100101",
    "01001100001101000100111000101111",
    "01001010001010111001000110100010",
    "01011101110010101101001010111000",
    "00110101000101010111010011000110",
    "11111001111100001100011011011110",
    "10111010000011111011001010111100",
    "11111101101100111010000110100001",
    "01011010011011100101110111010101",
    "01111110000111110100001101100010",
    "11000101101010000011000100011010",
    "11101100010000001100110010111100",
    "11000110101010101100111110011101",
    "10110110010010111101111110000011",
    "11111111010001110111011111100111",
    "11110110110000100001101111100100",
    "11010010110100010011010000101010",
    "10101011110101000011101111100100",
    "11100100110101011100001101101101",
    "10110000111000100100110100011111",
    "01000111011011110111111010111100",
    "11011100010011101001000000100011",
    "10101011111111110000010001000010",
    "10100001111101010101111000100001",
    "11111100110010010101010111101011",
    "01001100110000101011011011100110",
    "00110001000110100000100101111111",
    "01111110110001010001000000111001",
    "01001101110100100010000111101111",
    "01110010111110001000000110001000",
    "01010011000110100000011110110110",
    "00111100101101100011000110000001",
    "01100001011110100010011000010101",
    "11101110010111001100111100001011",
    "10111111101110011111010011001011",
    "10110001110000101001100000010010",
    "00001111100001100011010100010101",
    "01000011001111000000110101101001",
    "11010100010100100010100111110011",
    "01010010111110010000000000010010",
    "11111010000111100110101011000010",
    "01100010100100111100101001111110",
    "00010100100110110000001010011101",
    "01110011001100001100001011001000",
    "11011011110011010110011010100011",
    "10110011101100101101010010111001",
    "11011010000000010011110001001000",
    "01111010111001001000010100000010",
    "11010101100101010000001000010110",
    "01111001010010001101101010001000",
    "01000001001101011000011010101101",
    "11100001001000011100110101010100",
    "11010000110010100011011110100000",
    "11100000010110100101100011110110",
    "10100010010110010010011010011010",
    "01111101010001011010111100011010",
    "01111000001010011101010010100110",
    "01101110100010100101111010000011",
    "01011011000001010101010001101111",
    "11110011010000010111100000100101",
    "10110010110001000101011000011110",
    "01011011110100101101001000110101",
    "10011010011111111000001000010000",
    "11010101100101010100101000010010",
    "10110011110010001111101100010101",
    "01110101110000100110011100011010",
    "11011000001101101100101001000001");


  signal i : integer range 0 to n-1;
  signal j : std_logic;

  signal clk : std_logic;
  signal reset : std_logic;
  
  signal A, B, O : std_logic_vector(31 downto 0);

  signal count : integer range 0 to 3;
  
begin  -- STRUCTURE
  
  ibufg_inst : ibufg port map (I => clkin, O => clk);
  roc_inst : roc port map (O => reset);

  fa : FP_ADD port map (A => A, B => B, O => O);
  
  process (clk, reset)
  begin  -- process
    if reset = '1' then
      i <= 0;
      j <= '0';
      ledout <= "00";
    elsif clk'event and clk = '1' then
      if count = 0 then  
        -- count ��0�̎��̂ݎ��̍s�����s���i�N���b�N��1/4�{���Ɂj
        
        if j = '0' then
          -- j��0  ->  �o�͂���v���Ă��邩����
          if O /= table_o(i) then
            ledout(0) <= '1';
          end if;
          
          j <= '1';
        else
          -- j��1  ->  ���̃f�[�^��
          if i + 1 = n then
            i <= 0;
            ledout(1) <= '1';           -- �I���I
          else
            i <= i + 1;
          end if;

          j <= '0';
        end if;        
      end if;

      if count = 3 then
        count <= 0;
      else
        count <= count + 1;
      end if;
    end if;
    
    A <= table_a(i);
    B <= table_b(i);
  end process;
  
end STRUCTURE;
