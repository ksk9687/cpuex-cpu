library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

library unisim;
use unisim.vcomponents.all;

entity FP_CMP_TESTER is
  
  port (
    clkin  : in  std_logic;
    ledout : out std_logic);
    
end FP_CMP_TESTER;


architecture STRUCTURE of FP_CMP_TESTER is

  component FP_CMP
    port (
      A, B : in  std_logic_vector(31 downto 0);
      O    : out std_logic_vector(31 downto 0));
  end component;

  constant n : integer := 24;
  
  subtype vec32 is std_logic_vector(31 downto 0);
  type table32 is array(0 to n - 1) of vec32;
  
  constant table_a : table32 := (
    -- 0 vs 0
    "00000000000000000000000000000000",  -- +0.0
    "00000000000000000000000000000000",  -- +0.0
    "10000000000000000000000000000000",  -- -0.0
    "10000000000000000000000000000000",  -- -0.0

    -- 0 vs 1
    "00000000000000000000000000000000",  -- +0.0
    "00000000000000000000000000000000",  -- +0.0
    "10000000000000000000000000000000",  -- -0.0
    "10000000000000000000000000000000",  -- -0.0

    -- 1 vs 0
    "00111111100000000000000000000000",  -- +1.0
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0
    "10111111100000000000000000000000",  -- -1.0

    -- 1 vs 1
    "00111111100000000000000000000000",  -- +1.0
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0
    "10111111100000000000000000000000",  -- -1.0

    -- 1 vs 2
    "00111111100000000000000000000000",  -- +1.0
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0
    "10111111100000000000000000000000",  -- -1.0

    -- 2 vs 1
    "01000000000000000000000000000000",  -- +2.0
    "01000000000000000000000000000000",  -- +2.0
    "11000000000000000000000000000000",  -- -2.0
    "11000000000000000000000000000000"  -- -2.0
    );
  
  constant table_b : table32 := (
    -- 0 vs 0
    "00000000000000000000000000000000",  -- +0.0
    "10000000000000000000000000000000",  -- -0.0
    "00000000000000000000000000000000",  -- +0.0
    "10000000000000000000000000000000",  -- -0.0

    -- 0 vs 1
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0

    -- 1 vs 0
    "00000000000000000000000000000000",  -- +0.0
    "10000000000000000000000000000000",  -- -0.0
    "00000000000000000000000000000000",  -- +0.0
    "10000000000000000000000000000000",  -- -0.0

    -- 1 vs 1
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0

    -- 1 vs 2
    "01000000000000000000000000000000",  -- +2.0
    "11000000000000000000000000000000",  -- -2.0
    "01000000000000000000000000000000",  -- +2.0
    "11000000000000000000000000000000",  -- -2.0

    -- 2 vs 1
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000",  -- -1.0
    "00111111100000000000000000000000",  -- +1.0
    "10111111100000000000000000000000"  -- -1.0
    );
  
  signal clk, reset : std_logic;
  signal i : integer range 0 to n - 1;
  
  signal a, b, c : std_logic_vector(31 downto 0)
    := "00000000000000000000000000000000";
  
begin  -- STRUCTURE

  ibufg_inst : ibufg port map (I => clkin, O => clk);
  roc_inst : roc port map (O => reset);

  fp_cmp_inst : FP_CMP port map (A  => a, B  => b, O => c);

  ledout <= '0';

  process (clk, reset)
  begin  -- process
    if reset = '1' then
      i <= 0;

    elsif clk'event and clk = '1' then
      if i+1 = n then
        i <= 0;
      else
        i <= i+1;
      end if;
    end if;

    a <= table_a(i);
    b <= table_b(i);
  end process;
  
end STRUCTURE;
