library IEEE;
use IEEE.std_logic_1164.all;

library work;

package fp_sqrt_table is

subtype vec24 is std_logic_vector(23 downto 0);
type table_t is array (0 to 2047) of vec24;
constant table : table_t := (
"111111111111000000000001",
"111111111101000000001101",
"111111111011000000100101",
"111111111001000001001001",
"111111110111000001111001",
"111111110101000010110100",
"111111110011000011111100",
"111111110001000101001111",
"111111101111000110101110",
"111111101101001000011001",
"111111101011001010001111",
"111111101001001100010010",
"111111100111001110100000",
"111111100101010000111001",
"111111100011010011011110",
"111111100001010110001111",
"111111011111011001001011",
"111111011101011100010011",
"111111011011011111100111",
"111111011001100011000101",
"111111010111100110110000",
"111111010101101010100101",
"111111010011101110100110",
"111111010001110010110011",
"111111001111110111001011",
"111111001101111011101110",
"111111001100000000011100",
"111111001010000101010110",
"111111001000001010011011",
"111111000110001111101011",
"111111000100010101000110",
"111111000010011010101100",
"111111000000100000011110",
"111110111110100110011011",
"111110111100101100100010",
"111110111010110010110101",
"111110111000111001010011",
"111110110110111111111011",
"111110110101000110101111",
"111110110011001101101110",
"111110110001010100110111",
"111110101111011100001100",
"111110101101100011101011",
"111110101011101011010101",
"111110101001110011001010",
"111110100111111011001010",
"111110100110000011010101",
"111110100100001011101010",
"111110100010010100001010",
"111110100000011100110101",
"111110011110100101101010",
"111110011100101110101010",
"111110011010110111110101",
"111110011001000001001010",
"111110010111001010101010",
"111110010101010100010100",
"111110010011011110001001",
"111110010001101000001000",
"111110001111110010010010",
"111110001101111100100110",
"111110001100000111000101",
"111110001010010001101110",
"111110001000011100100001",
"111110000110100111011111",
"111110000100110010100111",
"111110000010111101111001",
"111110000001001001010110",
"111101111111010100111101",
"111101111101100000101110",
"111101111011101100101010",
"111101111001111000101111",
"111101111000000100111111",
"111101110110010001011001",
"111101110100011101111101",
"111101110010101010101011",
"111101110000110111100011",
"111101101111000100100101",
"111101101101010001110001",
"111101101011011111000111",
"111101101001101100100111",
"111101100111111010010001",
"111101100110001000000110",
"111101100100010110000011",
"111101100010100100001011",
"111101100000110010011101",
"111101011111000000111001",
"111101011101001111011110",
"111101011011011110001101",
"111101011001101101000110",
"111101010111111100001001",
"111101010110001011010101",
"111101010100011010101011",
"111101010010101010001011",
"111101010000111001110100",
"111101001111001001101000",
"111101001101011001100100",
"111101001011101001101011",
"111101001001111001111011",
"111101001000001010010100",
"111101000110011010110111",
"111101000100101011100100",
"111101000010111100011010",
"111101000001001101011001",
"111100111111011110100010",
"111100111101101111110101",
"111100111100000001010000",
"111100111010010010110110",
"111100111000100100100100",
"111100110110110110011100",
"111100110101001000011101",
"111100110011011010101000",
"111100110001101100111100",
"111100101111111111011001",
"111100101110010001111111",
"111100101100100100101111",
"111100101010110111101000",
"111100101001001010101010",
"111100100111011101110101",
"111100100101110001001001",
"111100100100000100100111",
"111100100010011000001101",
"111100100000101011111101",
"111100011110111111110101",
"111100011101010011110111",
"111100011011101000000010",
"111100011001111100010110",
"111100011000010000110010",
"111100010110100101011000",
"111100010100111010000111",
"111100010011001110111110",
"111100010001100011111111",
"111100001111111001001000",
"111100001110001110011011",
"111100001100100011110110",
"111100001010111001011010",
"111100001001001111000111",
"111100000111100100111100",
"111100000101111010111010",
"111100000100010001000010",
"111100000010100111010001",
"111100000000111101101010",
"111011111111010100001011",
"111011111101101010110101",
"111011111100000001101000",
"111011111010011000100011",
"111011111000101111100111",
"111011110111000110110011",
"111011110101011110001001",
"111011110011110101100110",
"111011110010001101001100",
"111011110000100100111011",
"111011101110111100110010",
"111011101101010100110010",
"111011101011101100111010",
"111011101010000101001011",
"111011101000011101100100",
"111011100110110110000110",
"111011100101001110110000",
"111011100011100111100010",
"111011100010000000011101",
"111011100000011001100000",
"111011011110110010101100",
"111011011101001011111111",
"111011011011100101011011",
"111011011001111111000000",
"111011011000011000101100",
"111011010110110010100001",
"111011010101001100011110",
"111011010011100110100100",
"111011010010000000110001",
"111011010000011011000111",
"111011001110110101100101",
"111011001101010000001011",
"111011001011101010111001",
"111011001010000101101111",
"111011001000100000101110",
"111011000110111011110100",
"111011000101010111000011",
"111011000011110010011001",
"111011000010001101111000",
"111011000000101001011110",
"111010111111000101001101",
"111010111101100001000011",
"111010111011111101000010",
"111010111010011001001000",
"111010111000110101010111",
"111010110111010001101101",
"111010110101101110001011",
"111010110100001010110010",
"111010110010100111100000",
"111010110001000100010101",
"111010101111100001010011",
"111010101101111110011000",
"111010101100011011100110",
"111010101010111000111011",
"111010101001010110011000",
"111010100111110011111100",
"111010100110010001101001",
"111010100100101111011101",
"111010100011001101011000",
"111010100001101011011100",
"111010100000001001100111",
"111010011110100111111010",
"111010011101000110010100",
"111010011011100100110110",
"111010011010000011100000",
"111010011000100010010001",
"111010010111000001001010",
"111010010101100000001010",
"111010010011111111010010",
"111010010010011110100010",
"111010010000111101111001",
"111010001111011101010111",
"111010001101111100111101",
"111010001100011100101011",
"111010001010111100100000",
"111010001001011100011100",
"111010000111111100100000",
"111010000110011100101011",
"111010000100111100111110",
"111010000011011101011000",
"111010000001111101111001",
"111010000000011110100010",
"111001111110111111010010",
"111001111101100000001001",
"111001111100000001001000",
"111001111010100010001110",
"111001111001000011011011",
"111001110111100100110000",
"111001110110000110001100",
"111001110100100111101111",
"111001110011001001011001",
"111001110001101011001010",
"111001110000001101000011",
"111001101110101111000011",
"111001101101010001001010",
"111001101011110011011000",
"111001101010010101101101",
"111001101000111000001010",
"111001100111011010101101",
"111001100101111101011000",
"111001100100100000001010",
"111001100011000011000010",
"111001100001100110000010",
"111001100000001001001001",
"111001011110101100010111",
"111001011101001111101100",
"111001011011110011001000",
"111001011010010110101011",
"111001011000111010010101",
"111001010111011110000101",
"111001010110000001111101",
"111001010100100101111100",
"111001010011001010000001",
"111001010001101110001110",
"111001010000010010100001",
"111001001110110110111100",
"111001001101011011011101",
"111001001100000000000101",
"111001001010100100110100",
"111001001001001001101001",
"111001000111101110100110",
"111001000110010011101001",
"111001000100111000110011",
"111001000011011110000100",
"111001000010000011011011",
"111001000000101000111010",
"111000111111001110011111",
"111000111101110100001011",
"111000111100011001111101",
"111000111010111111110110",
"111000111001100101110110",
"111000111000001011111100",
"111000110110110010001010",
"111000110101011000011101",
"111000110011111110111000",
"111000110010100101011001",
"111000110001001100000000",
"111000101111110010101111",
"111000101110011001100100",
"111000101101000000011111",
"111000101011100111100001",
"111000101010001110101001",
"111000101000110101111000",
"111000100111011101001110",
"111000100110000100101010",
"111000100100101100001100",
"111000100011010011110101",
"111000100001111011100101",
"111000100000100011011010",
"111000011111001011010111",
"111000011101110011011001",
"111000011100011011100011",
"111000011011000011110010",
"111000011001101100001000",
"111000011000010100100100",
"111000010110111101000111",
"111000010101100101110000",
"111000010100001110100000",
"111000010010110111010101",
"111000010001100000010001",
"111000010000001001010100",
"111000001110110010011100",
"111000001101011011101011",
"111000001100000101000000",
"111000001010101110011100",
"111000001001010111111110",
"111000001000000001100110",
"111000000110101011010100",
"111000000101010101001000",
"111000000011111111000011",
"111000000010101001000011",
"111000000001010011001010",
"110111111111111101011000",
"110111111110100111101011",
"110111111101010010000100",
"110111111011111100100100",
"110111111010100111001001",
"110111111001010001110101",
"110111110111111100100111",
"110111110110100111011111",
"110111110101010010011101",
"110111110011111101100001",
"110111110010101000101011",
"110111110001010011111011",
"110111101111111111010010",
"110111101110101010101110",
"110111101101010110010000",
"110111101100000001111000",
"110111101010101101100111",
"110111101001011001011011",
"110111101000000101010101",
"110111100110110001010101",
"110111100101011101011011",
"110111100100001001100111",
"110111100010110101111001",
"110111100001100010010001",
"110111100000001110101110",
"110111011110111011010010",
"110111011101100111111100",
"110111011100010100101011",
"110111011011000001100000",
"110111011001101110011011",
"110111011000011011011100",
"110111010111001000100011",
"110111010101110101101111",
"110111010100100011000001",
"110111010011010000011010",
"110111010001111101110111",
"110111010000101011011011",
"110111001111011001000100",
"110111001110000110110100",
"110111001100110100101000",
"110111001011100010100011",
"110111001010010000100011",
"110111001000111110101001",
"110111000111101100110101",
"110111000110011011000111",
"110111000101001001011110",
"110111000011110111111011",
"110111000010100110011101",
"110111000001010101000101",
"110111000000000011110011",
"110110111110110010100110",
"110110111101100001011111",
"110110111100010000011110",
"110110111010111111100010",
"110110111001101110101011",
"110110111000011101111011",
"110110110111001101010000",
"110110110101111100101010",
"110110110100101100001010",
"110110110011011011101111",
"110110110010001011011010",
"110110110000111011001011",
"110110101111101011000001",
"110110101110011010111101",
"110110101101001010111110",
"110110101011111011000100",
"110110101010101011010000",
"110110101001011011100010",
"110110101000001011111000",
"110110100110111100010101",
"110110100101101100110110",
"110110100100011101011110",
"110110100011001110001010",
"110110100001111110111100",
"110110100000101111110100",
"110110011111100000110000",
"110110011110010001110010",
"110110011101000010111010",
"110110011011110100000111",
"110110011010100101011001",
"110110011001010110110000",
"110110011000001000001101",
"110110010110111001101111",
"110110010101101011010111",
"110110010100011101000011",
"110110010011001110110101",
"110110010010000000101101",
"110110010000110010101001",
"110110001111100100101011",
"110110001110010110110010",
"110110001101001000111110",
"110110001011111011010000",
"110110001010101101100111",
"110110001001100000000011",
"110110001000010010100100",
"110110000111000101001010",
"110110000101110111110110",
"110110000100101010100110",
"110110000011011101011100",
"110110000010010000010111",
"110110000001000011010111",
"110101111111110110011101",
"110101111110101001100111",
"110101111101011100110111",
"110101111100010000001011",
"110101111011000011100101",
"110101111001110111000100",
"110101111000101010101000",
"110101110111011110010001",
"110101110110010001111111",
"110101110101000101110010",
"110101110011111001101011",
"110101110010101101101000",
"110101110001100001101010",
"110101110000010101110001",
"110101101111001001111110",
"110101101101111110001111",
"110101101100110010100110",
"110101101011100111000001",
"110101101010011011100001",
"110101101001010000000110",
"110101101000000100110001",
"110101100110111001100000",
"110101100101101110010100",
"110101100100100011001101",
"110101100011011000001011",
"110101100010001101001110",
"110101100001000010010110",
"110101011111110111100011",
"110101011110101100110101",
"110101011101100010001011",
"110101011100010111100111",
"110101011011001101000111",
"110101011010000010101100",
"110101011000111000010110",
"110101010111101110000101",
"110101010110100011111001",
"110101010101011001110001",
"110101010100001111101111",
"110101010011000101110001",
"110101010001111011111000",
"110101010000110010000100",
"110101001111101000010100",
"110101001110011110101010",
"110101001101010101000100",
"110101001100001011100011",
"110101001011000010000110",
"110101001001111000101111",
"110101001000101111011100",
"110101000111100110001110",
"110101000110011101000100",
"110101000101010100000000",
"110101000100001011000000",
"110101000011000010000101",
"110101000001111001001110",
"110101000000110000011100",
"110100111111100111101111",
"110100111110011111000111",
"110100111101010110100011",
"110100111100001110000011",
"110100111011000101101001",
"110100111001111101010011",
"110100111000110101000010",
"110100110111101100110101",
"110100110110100100101101",
"110100110101011100101010",
"110100110100010100101011",
"110100110011001100110001",
"110100110010000100111011",
"110100110000111101001010",
"110100101111110101011101",
"110100101110101101110101",
"110100101101100110010010",
"110100101100011110110011",
"110100101011010111011001",
"110100101010010000000011",
"110100101001001000110010",
"110100101000000001100101",
"110100100110111010011101",
"110100100101110011011001",
"110100100100101100011010",
"110100100011100101100000",
"110100100010011110101001",
"110100100001010111111000",
"110100100000010001001010",
"110100011111001010100001",
"110100011110000011111101",
"110100011100111101011101",
"110100011011110111000010",
"110100011010110000101011",
"110100011001101010011000",
"110100011000100100001010",
"110100010111011110000000",
"110100010110010111111010",
"110100010101010001111001",
"110100010100001011111101",
"110100010011000110000101",
"110100010010000000010001",
"110100010000111010100001",
"110100001111110100110110",
"110100001110101111001111",
"110100001101101001101101",
"110100001100100100001111",
"110100001011011110110101",
"110100001010011001011111",
"110100001001010100001110",
"110100001000001111000001",
"110100000111001001111001",
"110100000110000100110100",
"110100000100111111110101",
"110100000011111010111001",
"110100000010110110000001",
"110100000001110001001110",
"110100000000101100011111",
"110011111111100111110101",
"110011111110100011001110",
"110011111101011110101100",
"110011111100011010001110",
"110011111011010101110101",
"110011111010010001011111",
"110011111001001101001110",
"110011111000001001000001",
"110011110111000100111000",
"110011110110000000110011",
"110011110100111100110011",
"110011110011111000110111",
"110011110010110100111111",
"110011110001110001001011",
"110011110000101101011011",
"110011101111101001101111",
"110011101110100110001000",
"110011101101100010100100",
"110011101100011111000101",
"110011101011011011101010",
"110011101010011000010011",
"110011101001010101000000",
"110011101000010001110001",
"110011100111001110100111",
"110011100110001011100000",
"110011100101001000011110",
"110011100100000101011111",
"110011100011000010100101",
"110011100001111111101111",
"110011100000111100111101",
"110011011111111010001110",
"110011011110110111100100",
"110011011101110100111110",
"110011011100110010011100",
"110011011011101111111110",
"110011011010101101100100",
"110011011001101011001110",
"110011011000101000111100",
"110011010111100110101110",
"110011010110100100100101",
"110011010101100010011111",
"110011010100100000011101",
"110011010011011110011111",
"110011010010011100100101",
"110011010001011010101111",
"110011010000011000111100",
"110011001111010111001110",
"110011001110010101100100",
"110011001101010011111110",
"110011001100010010011100",
"110011001011010000111101",
"110011001010001111100011",
"110011001001001110001100",
"110011001000001100111010",
"110011000111001011101011",
"110011000110001010100000",
"110011000101001001011001",
"110011000100001000010110",
"110011000011000111010111",
"110011000010000110011100",
"110011000001000101100100",
"110011000000000100110001",
"110010111111000100000001",
"110010111110000011010101",
"110010111101000010101101",
"110010111100000010001001",
"110010111011000001101001",
"110010111010000001001100",
"110010111001000000110011",
"110010111000000000011111",
"110010110111000000001110",
"110010110110000000000000",
"110010110100111111110111",
"110010110011111111110001",
"110010110010111111101111",
"110010110001111111110001",
"110010110000111111110111",
"110010110000000000000000",
"110010101111000000001101",
"110010101110000000011110",
"110010101101000000110011",
"110010101100000001001100",
"110010101011000001101000",
"110010101010000010001000",
"110010101001000010101011",
"110010101000000011010011",
"110010100111000011111110",
"110010100110000100101101",
"110010100101000101011111",
"110010100100000110010101",
"110010100011000111001111",
"110010100010001000001101",
"110010100001001001001110",
"110010100000001010010011",
"110010011111001011011100",
"110010011110001100101000",
"110010011101001101111000",
"110010011100001111001011",
"110010011011010000100011",
"110010011010010001111110",
"110010011001010011011100",
"110010011000010100111110",
"110010010111010110100100",
"110010010110011000001110",
"110010010101011001111011",
"110010010100011011101011",
"110010010011011101011111",
"110010010010011111010111",
"110010010001100001010011",
"110010010000100011010010",
"110010001111100101010100",
"110010001110100111011011",
"110010001101101001100100",
"110010001100101011110010",
"110010001011101110000011",
"110010001010110000010111",
"110010001001110010101111",
"110010001000110101001011",
"110010000111110111101010",
"110010000110111010001100",
"110010000101111100110010",
"110010000100111111011100",
"110010000100000010001001",
"110010000011000100111010",
"110010000010000111101110",
"110010000001001010100110",
"110010000000001101100001",
"110001111111010000100000",
"110001111110010011100010",
"110001111101010110101000",
"110001111100011001110001",
"110001111011011100111110",
"110001111010100000001110",
"110001111001100011100001",
"110001111000100110111000",
"110001110111101010010011",
"110001110110101101110001",
"110001110101110001010010",
"110001110100110100110111",
"110001110011111000011111",
"110001110010111100001011",
"110001110001111111111010",
"110001110001000011101100",
"110001110000000111100010",
"110001101111001011011100",
"110001101110001111011000",
"110001101101010011011001",
"110001101100010111011100",
"110001101011011011100011",
"110001101010011111101101",
"110001101001100011111011",
"110001101000101000001100",
"110001100111101100100000",
"110001100110110000111000",
"110001100101110101010011",
"110001100100111001110010",
"110001100011111110010100",
"110001100011000010111001",
"110001100010000111100001",
"110001100001001100001101",
"110001100000010000111100",
"110001011111010101101111",
"110001011110011010100100",
"110001011101011111011110",
"110001011100100100011010",
"110001011011101001011010",
"110001011010101110011101",
"110001011001110011100011",
"110001011000111000101101",
"110001010111111101111010",
"110001010111000011001010",
"110001010110001000011101",
"110001010101001101110100",
"110001010100010011001110",
"110001010011011000101011",
"110001010010011110001100",
"110001010001100011101111",
"110001010000101001010110",
"110001001111101111000001",
"110001001110110100101110",
"110001001101111010011111",
"110001001101000000010011",
"110001001100000110001010",
"110001001011001100000100",
"110001001010010010000010",
"110001001001011000000011",
"110001001000011110000111",
"110001000111100100001110",
"110001000110101010011000",
"110001000101110000100110",
"110001000100110110110110",
"110001000011111101001010",
"110001000011000011100010",
"110001000010001001111100",
"110001000001010000011001",
"110001000000010110111010",
"110000111111011101011110",
"110000111110100100000101",
"110000111101101010101111",
"110000111100110001011100",
"110000111011111000001100",
"110000111010111111000000",
"110000111010000101110111",
"110000111001001100110000",
"110000111000010011101101",
"110000110111011010101101",
"110000110110100001110000",
"110000110101101000110111",
"110000110100110000000000",
"110000110011110111001100",
"110000110010111110011100",
"110000110010000101101111",
"110000110001001101000100",
"110000110000010100011101",
"110000101111011011111001",
"110000101110100011011000",
"110000101101101010111010",
"110000101100110010011111",
"110000101011111010000111",
"110000101011000001110010",
"110000101010001001100001",
"110000101001010001010010",
"110000101000011001000110",
"110000100111100000111110",
"110000100110101000111000",
"110000100101110000110110",
"110000100100111000110110",
"110000100100000000111010",
"110000100011001001000000",
"110000100010010001001010",
"110000100001011001010110",
"110000100000100001100110",
"110000011111101001111000",
"110000011110110010001110",
"110000011101111010100110",
"110000011101000011000010",
"110000011100001011100001",
"110000011011010100000010",
"110000011010011100100111",
"110000011001100101001110",
"110000011000101101111000",
"110000010111110110100110",
"110000010110111111010110",
"110000010110001000001001",
"110000010101010001000000",
"110000010100011001111001",
"110000010011100010110101",
"110000010010101011110100",
"110000010001110100110110",
"110000010000111101111011",
"110000010000000111000011",
"110000001111010000001110",
"110000001110011001011011",
"110000001101100010101100",
"110000001100101100000000",
"110000001011110101010110",
"110000001010111110101111",
"110000001010001000001100",
"110000001001010001101011",
"110000001000011011001101",
"110000000111100100110010",
"110000000110101110011010",
"110000000101111000000100",
"110000000101000001110010",
"110000000100001011100010",
"110000000011010101010110",
"110000000010011111001100",
"110000000001101001000101",
"110000000000110011000001",
"101111111111111101000000",
"101111111111000111000001",
"101111111110010001000110",
"101111111101011011001101",
"101111111100100101010111",
"101111111011101111100100",
"101111111010111001110100",
"101111111010000100000110",
"101111111001001110011100",
"101111111000011000110100",
"101111110111100011001111",
"101111110110101101101101",
"101111110101111000001101",
"101111110101000010110001",
"101111110100001101010111",
"101111110011011000000000",
"101111110010100010101100",
"101111110001101101011010",
"101111110000111000001100",
"101111110000000011000000",
"101111101111001101110111",
"101111101110011000110001",
"101111101101100011101101",
"101111101100101110101100",
"101111101011111001101110",
"101111101011000100110011",
"101111101010001111111011",
"101111101001011011000101",
"101111101000100110010010",
"101111100111110001100010",
"101111100110111100110100",
"101111100110001000001001",
"101111100101010011100001",
"101111100100011110111100",
"101111100011101010011001",
"101111100010110101111010",
"101111100010000001011100",
"101111100001001101000010",
"101111100000011000101010",
"101111011111100100010101",
"101111011110110000000011",
"101111011101111011110011",
"101111011101000111100110",
"101111011100010011011100",
"101111011011011111010100",
"101111011010101011010000",
"101111011001110111001101",
"101111011001000011001110",
"101111011000001111010001",
"101111010111011011010111",
"101111010110100111011111",
"101111010101110011101010",
"101111010100111111111000",
"101111010100001100001001",
"101111010011011000011100",
"101111010010100100110001",
"101111010001110001001010",
"101111010000111101100101",
"101111010000001010000010",
"101111001111010110100011",
"101111001110100011000110",
"101111001101101111101011",
"101111001100111100010011",
"101111001100001000111110",
"101111001011010101101011",
"101111001010100010011011",
"101111001001101111001110",
"101111001000111100000011",
"101111001000001000111011",
"101111000111010101110110",
"101111000110100010110011",
"101111000101101111110010",
"101111000100111100110100",
"101111000100001001111001",
"101111000011010111000000",
"101111000010100100001010",
"101111000001110001010111",
"101111000000111110100110",
"101111000000001011111000",
"101110111111011001001100",
"101110111110100110100011",
"101110111101110011111100",
"101110111101000001011000",
"101110111100001110110110",
"101110111011011100010111",
"101110111010101001111011",
"101110111001110111100001",
"101110111001000101001001",
"101110111000010010110101",
"101110110111100000100010",
"101110110110101110010010",
"101110110101111100000101",
"101110110101001001111010",
"101110110100010111110010",
"101110110011100101101100",
"101110110010110011101001",
"101110110010000001101001",
"101110110001001111101010",
"101110110000011101101111",
"101110101111101011110101",
"101110101110111001111111",
"101110101110001000001010",
"101110101101010110011001",
"101110101100100100101001",
"101110101011110010111101",
"101110101011000001010010",
"101110101010001111101011",
"101110101001011110000101",
"101110101000101100100010",
"101110100111111011000010",
"101110100111001001100100",
"101110100110011000001000",
"101110100101100110101111",
"101110100100110101011001",
"101110100100000100000101",
"101110100011010010110011",
"101110100010100001100100",
"101110100001110000010111",
"101110100000111111001101",
"101110100000001110000101",
"101110011111011100111111",
"101110011110101011111100",
"101110011101111010111011",
"101110011101001001111101",
"101110011100011001000001",
"101110011011101000001000",
"101110011010110111010001",
"101110011010000110011100",
"101110011001010101101010",
"101110011000100100111011",
"101110010111110100001101",
"101110010111000011100010",
"101110010110010010111010",
"101110010101100010010011",
"101110010100110001110000",
"101110010100000001001110",
"101110010011010000101111",
"101110010010100000010011",
"101110010001101111111000",
"101110010000111111100000",
"101110010000001111001011",
"101110001111011110111000",
"101110001110101110100111",
"101110001101111110011000",
"101110001101001110001100",
"101110001100011110000011",
"101110001011101101111011",
"101110001010111101110110",
"101110001010001101110011",
"101110001001011101110011",
"101110001000101101110101",
"101110000111111101111001",
"101110000111001110000000",
"101110000110011110001001",
"101110000101101110010100",
"101110000100111110100010",
"101110000100001110110010",
"101110000011011111000100",
"101110000010101111011001",
"101110000001111111110000",
"101110000001010000001001",
"101110000000100000100100",
"101101111111110001000010",
"101101111111000001100010",
"101101111110010010000101",
"101101111101100010101010",
"101101111100110011010001",
"101101111100000011111010",
"101101111011010100100101",
"101101111010100101010011",
"101101111001110110000011",
"101101111001000110110110",
"101101111000010111101011",
"101101110111101000100010",
"101101110110111001011011",
"101101110110001010010110",
"101101110101011011010100",
"101101110100101100010100",
"101101110011111101010110",
"101101110011001110011011",
"101101110010011111100010",
"101101110001110000101011",
"101101110001000001110110",
"101101110000010011000100",
"101101101111100100010011",
"101101101110110101100101",
"101101101110000110111010",
"101101101101011000010000",
"101101101100101001101001",
"101101101011111011000100",
"101101101011001100100001",
"101101101010011110000000",
"101101101001101111100010",
"101101101001000001000110",
"101101101000010010101100",
"101101100111100100010100",
"101101100110110101111111",
"101101100110000111101011",
"101101100101011001011010",
"101101100100101011001011",
"101101100011111100111110",
"101101100011001110110100",
"101101100010100000101100",
"101101100001110010100101",
"101101100001000100100001",
"101101100000010110100000",
"101101011111101000100000",
"101101011110111010100011",
"101101011110001100100111",
"101101011101011110101110",
"101101011100110000110111",
"101101011100000011000011",
"101101011011010101010000",
"101101011010100111100000",
"101101011001111001110001",
"101101011001001100000101",
"101101011000011110011011",
"101101010111110000110011",
"101101010111000011001110",
"101101010110010101101010",
"101101010101101000001001",
"101101010100111010101010",
"101101010100001101001101",
"101101010011011111110010",
"101101010010110010011001",
"101101010010000101000010",
"101101010001010111101110",
"101101010000101010011011",
"101101001111100110100011",
"101101001110001100001011",
"101101001100110001111100",
"101101001011010111110100",
"101101001001111101110110",
"101101001000100011111111",
"101101000111001010010001",
"101101000101110000101011",
"101101000100010111001110",
"101101000010111101111001",
"101101000001100100101100",
"101101000000001011100111",
"101100111110110010101011",
"101100111101011001110111",
"101100111100000001001011",
"101100111010101000101000",
"101100111001010000001100",
"101100110111110111111001",
"101100110110011111101110",
"101100110101000111101011",
"101100110011101111110000",
"101100110010010111111101",
"101100110001000000010010",
"101100101111101000101111",
"101100101110010001010100",
"101100101100111010000010",
"101100101011100010110111",
"101100101010001011110100",
"101100101000110100111001",
"101100100111011110000110",
"101100100110000111011011",
"101100100100110000111000",
"101100100011011010011101",
"101100100010000100001001",
"101100100000101101111101",
"101100011111010111111010",
"101100011110000001111110",
"101100011100101100001001",
"101100011011010110011101",
"101100011010000000111000",
"101100011000101011011011",
"101100010111010110000110",
"101100010110000000111000",
"101100010100101011110010",
"101100010011010110110100",
"101100010010000001111101",
"101100010000101101001110",
"101100001111011000100110",
"101100001110000100000110",
"101100001100101111101110",
"101100001011011011011101",
"101100001010000111010100",
"101100001000110011010010",
"101100000111011111010111",
"101100000110001011100101",
"101100000100110111111001",
"101100000011100100010101",
"101100000010010000111001",
"101100000000111101100100",
"101011111111101010010110",
"101011111110010111001111",
"101011111101000100010000",
"101011111011110001011001",
"101011111010011110101000",
"101011111001001011111111",
"101011110111111001011101",
"101011110110100111000011",
"101011110101010100101111",
"101011110100000010100011",
"101011110010110000011111",
"101011110001011110100001",
"101011110000001100101010",
"101011101110111010111011",
"101011101101101001010011",
"101011101100010111110010",
"101011101011000110011000",
"101011101001110101000101",
"101011101000100011111010",
"101011100111010010110101",
"101011100110000001110111",
"101011100100110001000001",
"101011100011100000010001",
"101011100010001111101001",
"101011100000111111000111",
"101011011111101110101101",
"101011011110011110011001",
"101011011101001110001101",
"101011011011111110000111",
"101011011010101110001000",
"101011011001011110010000",
"101011011000001110011111",
"101011010110111110110101",
"101011010101101111010010",
"101011010100011111110101",
"101011010011010000100000",
"101011010010000001010001",
"101011010000110010001001",
"101011001111100011000111",
"101011001110010100001101",
"101011001101000101011001",
"101011001011110110101100",
"101011001010101000000110",
"101011001001011001100110",
"101011001000001011001101",
"101011000110111100111011",
"101011000101101110101111",
"101011000100100000101010",
"101011000011010010101100",
"101011000010000100110100",
"101011000000110111000011",
"101010111111101001011001",
"101010111110011011110101",
"101010111101001110010111",
"101010111100000001000000",
"101010111010110011110000",
"101010111001100110100110",
"101010111000011001100011",
"101010110111001100100110",
"101010110101111111101111",
"101010110100110010111111",
"101010110011100110010110",
"101010110010011001110011",
"101010110001001101010110",
"101010110000000001000000",
"101010101110110100110000",
"101010101101101000100110",
"101010101100011100100011",
"101010101011010000100110",
"101010101010000100110000",
"101010101000111000111111",
"101010100111101101010110",
"101010100110100001110010",
"101010100101010110010101",
"101010100100001010111110",
"101010100010111111101101",
"101010100001110100100010",
"101010100000101001011110",
"101010011111011110100000",
"101010011110010011101000",
"101010011101001000110110",
"101010011011111110001010",
"101010011010110011100101",
"101010011001101001000101",
"101010011000011110101100",
"101010010111010100011001",
"101010010110001010001100",
"101010010101000000000101",
"101010010011110110000100",
"101010010010101100001001",
"101010010001100010010101",
"101010010000011000100110",
"101010001111001110111101",
"101010001110000101011011",
"101010001100111011111110",
"101010001011110010100111",
"101010001010101001010110",
"101010001001100000001100",
"101010001000010111000111",
"101010000111001110001000",
"101010000110000101001111",
"101010000100111100011100",
"101010000011110011101111",
"101010000010101011001000",
"101010000001100010100110",
"101010000000011010001011",
"101001111111010001110101",
"101001111110001001100101",
"101001111101000001011011",
"101001111011111001010111",
"101001111010110001011000",
"101001111001101001100000",
"101001111000100001101101",
"101001110111011010000000",
"101001110110010010011000",
"101001110101001010110111",
"101001110100000011011011",
"101001110010111100000101",
"101001110001110100110100",
"101001110000101101101001",
"101001101111100110100100",
"101001101110011111100101",
"101001101101011000101011",
"101001101100010001110111",
"101001101011001011001000",
"101001101010000100100000",
"101001101000111101111100",
"101001100111110111011111",
"101001100110110001000110",
"101001100101101010110100",
"101001100100100100100111",
"101001100011011110100000",
"101001100010011000011110",
"101001100001010010100001",
"101001100000001100101010",
"101001011111000110111001",
"101001011110000001001101",
"101001011100111011100111",
"101001011011110110000110",
"101001011010110000101011",
"101001011001101011010101",
"101001011000100110000100",
"101001010111100000111001",
"101001010110011011110011",
"101001010101010110110011",
"101001010100010001111000",
"101001010011001101000011",
"101001010010001000010010",
"101001010001000011101000",
"101001001111111111000010",
"101001001110111010100010",
"101001001101110110000111",
"101001001100110001110010",
"101001001011101101100010",
"101001001010101001010111",
"101001001001100101010001",
"101001001000100001010001",
"101001000111011101010110",
"101001000110011001100000",
"101001000101010101110000",
"101001000100010010000100",
"101001000011001110011110",
"101001000010001010111101",
"101001000001000111100010",
"101001000000000100001011",
"101000111111000000111010",
"101000111101111101101110",
"101000111100111010100111",
"101000111011110111100101",
"101000111010110100101000",
"101000111001110001110001",
"101000111000101110111110",
"101000110111101100010001",
"101000110110101001101001",
"101000110101100111000110",
"101000110100100100101000",
"101000110011100010001111",
"101000110010011111111011",
"101000110001011101101100",
"101000110000011011100010",
"101000101111011001011101",
"101000101110010111011101",
"101000101101010101100011",
"101000101100010011101101",
"101000101011010001111100",
"101000101010010000010000",
"101000101001001110101001",
"101000101000001101000111",
"101000100111001011101010",
"101000100110001010010010",
"101000100101001000111111",
"101000100100000111110001",
"101000100011000110101000",
"101000100010000101100011",
"101000100001000100100100",
"101000100000000011101001",
"101000011111000010110100",
"101000011110000010000011",
"101000011101000001010111",
"101000011100000000110000",
"101000011011000000001101",
"101000011001111111110000",
"101000011000111111010111",
"101000010111111111000011",
"101000010110111110110100",
"101000010101111110101010",
"101000010100111110100100",
"101000010011111110100011",
"101000010010111110100111",
"101000010001111110110000",
"101000010000111110111110",
"101000001111111111010000",
"101000001110111111100111",
"101000001110000000000011",
"101000001101000000100011",
"101000001100000001001000",
"101000001011000001110010",
"101000001010000010100000",
"101000001001000011010011",
"101000001000000100001011",
"101000000111000101000111",
"101000000110000110001000",
"101000000101000111001110",
"101000000100001000011000",
"101000000011001001100111",
"101000000010001010111011",
"101000000001001100010011",
"101000000000001101110000",
"100111111111001111010001",
"100111111110010000110111",
"100111111101010010100001",
"100111111100010100010000",
"100111111011010110000100",
"100111111010010111111100",
"100111111001011001111000",
"100111111000011011111001",
"100111110111011101111111",
"100111110110100000001001",
"100111110101100010011000",
"100111110100100100101011",
"100111110011100111000010",
"100111110010101001011110",
"100111110001101011111111",
"100111110000101110100100",
"100111101111110001001101",
"100111101110110011111011",
"100111101101110110101101",
"100111101100111001100100",
"100111101011111100011111",
"100111101010111111011110",
"100111101010000010100010",
"100111101001000101101011",
"100111101000001000110111",
"100111100111001100001000",
"100111100110001111011110",
"100111100101010010110111",
"100111100100010110010101",
"100111100011011001111000",
"100111100010011101011110",
"100111100001100001001001",
"100111100000100100111001",
"100111011111101000101100",
"100111011110101100100100",
"100111011101110000100001",
"100111011100110100100001",
"100111011011111000100110",
"100111011010111100101111",
"100111011010000000111100",
"100111011001000101001110",
"100111011000001001100100",
"100111010111001101111110",
"100111010110010010011100",
"100111010101010110111110",
"100111010100011011100101",
"100111010011100000010000",
"100111010010100100111111",
"100111010001101001110010",
"100111010000101110101010",
"100111001111110011100101",
"100111001110111000100101",
"100111001101111101101001",
"100111001101000010110001",
"100111001100000111111101",
"100111001011001101001101",
"100111001010010010100010",
"100111001001010111111010",
"100111001000011101010111",
"100111000111100010111000",
"100111000110101000011101",
"100111000101101110000110",
"100111000100110011110011",
"100111000011111001100100",
"100111000010111111011001",
"100111000010000101010010",
"100111000001001011010000",
"100111000000010001010001",
"100110111111010111010110",
"100110111110011101100000",
"100110111101100011101101",
"100110111100101001111111",
"100110111011110000010100",
"100110111010110110101110",
"100110111001111101001011",
"100110111001000011101100",
"100110111000001010010010",
"100110110111010000111011",
"100110110110010111101001",
"100110110101011110011010",
"100110110100100101001111",
"100110110011101100001000",
"100110110010110011000101",
"100110110001111010000110",
"100110110001000001001011",
"100110110000001000010100",
"100110101111001111100001",
"100110101110010110110010",
"100110101101011110000110",
"100110101100100101011111",
"100110101011101100111011",
"100110101010110100011011",
"100110101001111011111111",
"100110101001000011100111",
"100110101000001011010011",
"100110100111010011000011",
"100110100110011010110110",
"100110100101100010101110",
"100110100100101010101001",
"100110100011110010101000",
"100110100010111010101010",
"100110100010000010110001",
"100110100001001010111011",
"100110100000010011001001",
"100110011111011011011011",
"100110011110100011110001",
"100110011101101100001011",
"100110011100110100101000",
"100110011011111101001001",
"100110011011000101101101",
"100110011010001110010110",
"100110011001010111000010",
"100110011000011111110010",
"100110010111101000100110",
"100110010110110001011101",
"100110010101111010011000",
"100110010101000011010111",
"100110010100001100011010",
"100110010011010101100000",
"100110010010011110101010",
"100110010001100111110111",
"100110010000110001001001",
"100110001111111010011101",
"100110001111000011110110",
"100110001110001101010010",
"100110001101010110110010",
"100110001100100000010110",
"100110001011101001111101",
"100110001010110011101000",
"100110001001111101010110",
"100110001001000111001000",
"100110001000010000111110",
"100110000111011010110111",
"100110000110100100110100",
"100110000101101110110100",
"100110000100111000111000",
"100110000100000011000000",
"100110000011001101001011",
"100110000010010111011001",
"100110000001100001101100",
"100110000000101100000001",
"100101111111110110011011",
"100101111111000000111000",
"100101111110001011011000",
"100101111101010101111100",
"100101111100100000100100",
"100101111011101011001111",
"100101111010110101111101",
"100101111010000000101111",
"100101111001001011100101",
"100101111000010110011110",
"100101110111100001011010",
"100101110110101100011010",
"100101110101110111011110",
"100101110101000010100101",
"100101110100001101101111",
"100101110011011000111101",
"100101110010100100001110",
"100101110001101111100011",
"100101110000111010111011",
"100101110000000110010111",
"100101101111010001110110",
"100101101110011101011000",
"100101101101101000111110",
"100101101100110100100111",
"100101101100000000010100",
"100101101011001100000100",
"100101101010010111111000",
"100101101001100011101110",
"100101101000101111101001",
"100101100111111011100110",
"100101100111000111100111",
"100101100110010011101100",
"100101100101011111110011",
"100101100100101011111110",
"100101100011111000001101",
"100101100011000100011111",
"100101100010010000110100",
"100101100001011101001100",
"100101100000101001101000",
"100101011111110110000111",
"100101011111000010101001",
"100101011110001111001111",
"100101011101011011111000",
"100101011100101000100100",
"100101011011110101010100",
"100101011011000010000111",
"100101011010001110111101",
"100101011001011011110111",
"100101011000101000110011",
"100101010111110101110011",
"100101010111000010110110",
"100101010110001111111101",
"100101010101011101000111",
"100101010100101010010100",
"100101010011110111100100",
"100101010011000100110111",
"100101010010010010001110",
"100101010001011111101000",
"100101010000101101000101",
"100101001111111010100101",
"100101001111001000001001",
"100101001110010101110000",
"100101001101100011011001",
"100101001100110001000111",
"100101001011111110110111",
"100101001011001100101010",
"100101001010011010100001",
"100101001001101000011011",
"100101001000110110011000",
"100101001000000100011000",
"100101000111010010011011",
"100101000110100000100010",
"100101000101101110101011",
"100101000100111100111000",
"100101000100001011001000",
"100101000011011001011011",
"100101000010100111110001",
"100101000001110110001010",
"100101000001000100100110",
"100101000000010011000110",
"100100111111100001101000",
"100100111110110000001110",
"100100111101111110110111",
"100100111101001101100011",
"100100111100011100010010",
"100100111011101011000011",
"100100111010111001111001",
"100100111010001000110001",
"100100111001010111101100",
"100100111000100110101010",
"100100110111110101101011",
"100100110111000100110000",
"100100110110010011110111",
"100100110101100011000001",
"100100110100110010001111",
"100100110100000001011111",
"100100110011010000110011",
"100100110010100000001001",
"100100110001101111100011",
"100100110000111110111111",
"100100110000001110011111",
"100100101111011110000001",
"100100101110101101100111",
"100100101101111101001111",
"100100101101001100111011",
"100100101100011100101001",
"100100101011101100011011",
"100100101010111100001111",
"100100101010001100000111",
"100100101001011100000001",
"100100101000101011111110",
"100100100111111011111111",
"100100100111001100000010",
"100100100110011100001000",
"100100100101101100010001",
"100100100100111100011101",
"100100100100001100101100",
"100100100011011100111110",
"100100100010101101010011",
"100100100001111101101010",
"100100100001001110000101",
"100100100000011110100010",
"100100011111101111000011",
"100100011110111111100110",
"100100011110010000001100",
"100100011101100000110101",
"100100011100110001100001",
"100100011100000010010000",
"100100011011010011000010",
"100100011010100011110110",
"100100011001110100101110",
"100100011001000101101000",
"100100011000010110100101",
"100100010111100111100101",
"100100010110111000101000",
"100100010110001001101101",
"100100010101011010110110",
"100100010100101100000001",
"100100010011111101001111",
"100100010011001110100000",
"100100010010011111110100",
"100100010001110001001011",
"100100010001000010100100",
"100100010000010100000000",
"100100001111100101011111",
"100100001110110111000001",
"100100001110001000100110",
"100100001101011010001101",
"100100001100101011110111",
"100100001011111101100100",
"100100001011001111010100",
"100100001010100001000111",
"100100001001110010111100",
"100100001001000100110100",
"100100001000010110101111",
"100100000111101000101100",
"100100000110111010101101",
"100100000110001100110000",
"100100000101011110110101",
"100100000100110000111110",
"100100000100000011001001",
"100100000011010101010111",
"100100000010100111101000",
"100100000001111001111011",
"100100000001001100010001",
"100100000000011110101010",
"100011111111110001000110",
"100011111111000011100100",
"100011111110010110000101",
"100011111101101000101000",
"100011111100111011001111",
"100011111100001101111000",
"100011111011100000100011",
"100011111010110011010010",
"100011111010000110000011",
"100011111001011000110111",
"100011111000101011101101",
"100011110111111110100110",
"100011110111010001100010",
"100011110110100100100000",
"100011110101110111100001",
"100011110101001010100101",
"100011110100011101101011",
"100011110011110000110100",
"100011110011000011111111",
"100011110010010111001101",
"100011110001101010011110",
"100011110000111101110010",
"100011110000010001001000",
"100011101111100100100000",
"100011101110110111111011",
"100011101110001011011001",
"100011101101011110111010",
"100011101100110010011101",
"100011101100000110000010",
"100011101011011001101011",
"100011101010101101010101",
"100011101010000001000011",
"100011101001010100110011",
"100011101000101000100101",
"100011100111111100011010",
"100011100111010000010010",
"100011100110100100001100",
"100011100101111000001001",
"100011100101001100001000",
"100011100100100000001010",
"100011100011110100001111",
"100011100011001000010110",
"100011100010011100011111",
"100011100001110000101011",
"100011100001000100111010",
"100011100000011001001011",
"100011011111101101011111",
"100011011111000001110101",
"100011011110010110001101",
"100011011101101010101001",
"100011011100111111000110",
"100011011100010011100110",
"100011011011101000001001",
"100011011010111100101110",
"100011011010010001010110",
"100011011001100110000000",
"100011011000111010101101",
"100011011000001111011100",
"100011010111100100001110",
"100011010110111001000010",
"100011010110001101111000",
"100011010101100010110001",
"100011010100110111101101",
"100011010100001100101011",
"100011010011100001101011",
"100011010010110110101110",
"100011010010001011110011",
"100011010001100000111011",
"100011010000110110000101",
"100011010000001011010010",
"100011001111100000100001",
"100011001110110101110010",
"100011001110001011000110",
"100011001101100000011101",
"100011001100110101110101",
"100011001100001011010000",
"100011001011100000101110",
"100011001010110110001110",
"100011001010001011110000",
"100011001001100001010101",
"100011001000110110111100",
"100011001000001100100110",
"100011000111100010010010",
"100011000110111000000000",
"100011000110001101110001",
"100011000101100011100100",
"100011000100111001011010",
"100011000100001111010010",
"100011000011100101001100",
"100011000010111011001001",
"100011000010010001000111",
"100011000001100111001001",
"100011000000111101001101",
"100011000000010011010011",
"100010111111101001011011",
"100010111110111111100110",
"100010111110010101110011",
"100010111101101100000010",
"100010111101000010010100",
"100010111100011000101000",
"100010111011101110111111",
"100010111011000101010111",
"100010111010011011110010",
"100010111001110010010000",
"100010111001001000110000",
"100010111000011111010010",
"100010110111110101110110",
"100010110111001100011101",
"100010110110100011000101",
"100010110101111001110001",
"100010110101010000011110",
"100010110100100111001110",
"100010110011111110000000",
"100010110011010100110101",
"100010110010101011101011",
"100010110010000010100100",
"100010110001011001011111",
"100010110000110000011101",
"100010110000000111011101",
"100010101111011110011111",
"100010101110110101100011",
"100010101110001100101010",
"100010101101100011110010",
"100010101100111010111110",
"100010101100010010001011",
"100010101011101001011010",
"100010101011000000101100",
"100010101010011000000000",
"100010101001101111010111",
"100010101001000110101111",
"100010101000011110001010",
"100010100111110101100111",
"100010100111001101000110",
"100010100110100100101000",
"100010100101111100001011",
"100010100101010011110001",
"100010100100101011011001",
"100010100100000011000011",
"100010100011011010110000",
"100010100010110010011111",
"100010100010001010001111",
"100010100001100010000011",
"100010100000111001111000",
"100010100000010001101111",
"100010011111101001101001",
"100010011111000001100101",
"100010011110011001100011",
"100010011101110001100011",
"100010011101001001100101",
"100010011100100001101010",
"100010011011111001110001",
"100010011011010001111001",
"100010011010101010000100",
"100010011010000010010010",
"100010011001011010100001",
"100010011000110010110010",
"100010011000001011000110",
"100010010111100011011100",
"100010010110111011110100",
"100010010110010100001110",
"100010010101101100101010",
"100010010101000101001000",
"100010010100011101101001",
"100010010011110110001100",
"100010010011001110110000",
"100010010010100111010111",
"100010010010000000000000",
"100010010001011000101011",
"100010010000110001011000",
"100010010000001010001000",
"100010001111100010111001",
"100010001110111011101101",
"100010001110010100100010",
"100010001101101101011010",
"100010001101000110010100",
"100010001100011111010000",
"100010001011111000001110",
"100010001011010001001110",
"100010001010101010010000",
"100010001010000011010100",
"100010001001011100011011",
"100010001000110101100011",
"100010001000001110101110",
"100010000111100111111010",
"100010000111000001001001",
"100010000110011010011001",
"100010000101110011101100",
"100010000101001101000001",
"100010000100100110011000",
"100010000011111111110001",
"100010000011011001001100",
"100010000010110010101001",
"100010000010001100001000",
"100010000001100101101001",
"100010000000111111001100",
"100010000000011000110001",
"100001111111110010011000",
"100001111111001100000010",
"100001111110100101101101",
"100001111101111111011010",
"100001111101011001001001",
"100001111100110010111011",
"100001111100001100101110",
"100001111011100110100011",
"100001111011000000011011",
"100001111010011010010100",
"100001111001110100010000",
"100001111001001110001101",
"100001111000101000001100",
"100001111000000010001110",
"100001110111011100010001",
"100001110110110110010111",
"100001110110010000011110",
"100001110101101010100111",
"100001110101000100110011",
"100001110100011111000000",
"100001110011111001001111",
"100001110011010011100000",
"100001110010101101110100",
"100001110010001000001001",
"100001110001100010100000",
"100001110000111100111001",
"100001110000010111010100",
"100001101111110001110001",
"100001101111001100010000",
"100001101110100110110001",
"100001101110000001010100",
"100001101101011011111001",
"100001101100110110100000",
"100001101100010001001001",
"100001101011101011110011",
"100001101011000110100000",
"100001101010100001001110",
"100001101001111011111111",
"100001101001010110110001",
"100001101000110001100110",
"100001101000001100011100",
"100001100111100111010100",
"100001100111000010001110",
"100001100110011101001010",
"100001100101111000001000",
"100001100101010011001000",
"100001100100101110001010",
"100001100100001001001110",
"100001100011100100010011",
"100001100010111111011011",
"100001100010011010100100",
"100001100001110101101111",
"100001100001010000111101",
"100001100000101100001100",
"100001100000000111011101",
"100001011111100010110000",
"100001011110111110000100",
"100001011110011001011011",
"100001011101110100110011",
"100001011101010000001110",
"100001011100101011101010",
"100001011100000111001000",
"100001011011100010101000",
"100001011010111110001010",
"100001011010011001101110",
"100001011001110101010011",
"100001011001010000111011",
"100001011000101100100100",
"100001011000001000001111",
"100001010111100011111100",
"100001010110111111101011",
"100001010110011011011100",
"100001010101110111001110",
"100001010101010011000011",
"100001010100101110111001",
"100001010100001010110001",
"100001010011100110101011",
"100001010011000010100110",
"100001010010011110100100",
"100001010001111010100011",
"100001010001010110100101",
"100001010000110010101000",
"100001010000001110101100",
"100001001111101010110011",
"100001001111000110111100",
"100001001110100011000110",
"100001001101111111010010",
"100001001101011011100000",
"100001001100110111110000",
"100001001100010100000001",
"100001001011110000010100",
"100001001011001100101010",
"100001001010101001000001",
"100001001010000101011001",
"100001001001100001110100",
"100001001000111110010000",
"100001001000011010101110",
"100001000111110111001110",
"100001000111010011110000",
"100001000110110000010011",
"100001000110001100111000",
"100001000101101001011111",
"100001000101000110001000",
"100001000100100010110011",
"100001000011111111011111",
"100001000011011100001101",
"100001000010111000111101",
"100001000010010101101110",
"100001000001110010100010",
"100001000001001111010111",
"100001000000101100001110",
"100001000000001001000110",
"100000111111100110000001",
"100000111111000010111101",
"100000111110011111111011",
"100000111101111100111010",
"100000111101011001111011",
"100000111100110110111111",
"100000111100010100000011",
"100000111011110001001010",
"100000111011001110010010",
"100000111010101011011100",
"100000111010001000101000",
"100000111001100101110101",
"100000111001000011000101",
"100000111000100000010101",
"100000110111111101101000",
"100000110111011010111100",
"100000110110111000010010",
"100000110110010101101010",
"100000110101110011000100",
"100000110101010000011111",
"100000110100101101111100",
"100000110100001011011010",
"100000110011101000111011",
"100000110011000110011101",
"100000110010100100000000",
"100000110010000001100110",
"100000110001011111001101",
"100000110000111100110110",
"100000110000011010100000",
"100000101111111000001100",
"100000101111010101111010",
"100000101110110011101001",
"100000101110010001011011",
"100000101101101111001110",
"100000101101001101000010",
"100000101100101010111000",
"100000101100001000110000",
"100000101011100110101010",
"100000101011000100100101",
"100000101010100010100010",
"100000101010000000100000",
"100000101001011110100001",
"100000101000111100100010",
"100000101000011010100110",
"100000100111111000101011",
"100000100111010110110010",
"100000100110110100111010",
"100000100110010011000101",
"100000100101110001010000",
"100000100101001111011110",
"100000100100101101101101",
"100000100100001011111101",
"100000100011101010010000",
"100000100011001000100100",
"100000100010100110111001",
"100000100010000101010001",
"100000100001100011101001",
"100000100001000010000100",
"100000100000100000100000",
"100000011111111110111110",
"100000011111011101011101",
"100000011110111011111110",
"100000011110011010100001",
"100000011101111001000101",
"100000011101010111101011",
"100000011100110110010010",
"100000011100010100111011",
"100000011011110011100110",
"100000011011010010010010",
"100000011010110001000000",
"100000011010001111101111",
"100000011001101110100000",
"100000011001001101010011",
"100000011000101100000111",
"100000011000001010111101",
"100000010111101001110100",
"100000010111001000101110",
"100000010110100111101000",
"100000010110000110100100",
"100000010101100101100010",
"100000010101000100100001",
"100000010100100011100010",
"100000010100000010100101",
"100000010011100001101001",
"100000010011000000101111",
"100000010010011111110110",
"100000010001111110111111",
"100000010001011110001001",
"100000010000111101010101",
"100000010000011100100010",
"100000001111111011110001",
"100000001111011011000010",
"100000001110111010010100",
"100000001110011001101000",
"100000001101111000111101",
"100000001101011000010100",
"100000001100110111101100",
"100000001100010111000110",
"100000001011110110100010",
"100000001011010101111111",
"100000001010110101011101",
"100000001010010100111101",
"100000001001110100011111",
"100000001001010100000010",
"100000001000110011100111",
"100000001000010011001101",
"100000000111110010110101",
"100000000111010010011110",
"100000000110110010001001",
"100000000110010001110101",
"100000000101110001100011",
"100000000101010001010011",
"100000000100110001000011",
"100000000100010000110110",
"100000000011110000101010",
"100000000011010000011111",
"100000000010110000010110",
"100000000010010000001111",
"100000000001110000001001",
"100000000001010000000100",
"100000000000110000000001",
"100000000000010000000000"
);

end package fp_sqrt_table;
